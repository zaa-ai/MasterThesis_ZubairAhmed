virtual clk_reset_if vif_clk_rst;

buffer_reader_action_e	action;

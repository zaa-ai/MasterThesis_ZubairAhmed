/* ###   interface instances   ###################################################### */

scan_registers_SCAN_if scan_registers_SCAN (); 


real TRIM__I5U__ = 0;
real TRIM__OT__ = 3;
real TRIM__DSI1_rx1_rise__ = 8;
real TRIM__DSI1_rx1_fall__ = 9;
real TRIM__DSI1_rx2_rise__ = 1;
real TRIM__DSI1_rx2_fall__ = 0;
real TRIM__DSI0_rx1_rise__ = 8;
real TRIM__DSI0_rx1_fall__ = 9;
real TRIM__DSI0_rx2_rise__ = 1;
real TRIM__DSI0_rx2_fall__ = 0;
real TRIM__OSC_F__ = 73;

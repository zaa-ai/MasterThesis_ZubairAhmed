
slave_timing[3][0].info_corner          = 1;
slave_timing[3][0].info_temp__j__       = 125;
slave_timing[3][0].info_i__quite_rec__  = 0.006000000;
slave_timing[3][0].info_dtr__ib__       = -1;
slave_timing[3][0].info_i__offset_rec__ = 0.000000000;
slave_timing[3][0].info_i__max_slave__  = 0.023000000;
slave_timing[3][0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][0].info_r__dsi_bus__    = 5.000;

slave_timing[3][0].t_rxd1[0][1] = 2745ns;
slave_timing[3][0].t_rxd1[1][0] = 2734ns;
slave_timing[3][0].t_rxd1[0][2] = 2054ns;
slave_timing[3][0].t_rxd1[2][0] = 3321ns;
slave_timing[3][0].t_rxd2[0][2] = 3289ns;
slave_timing[3][0].t_rxd2[2][0] = 2032ns;
slave_timing[3][0].t_rxd2[1][2] = 2720ns;
slave_timing[3][0].t_rxd2[2][1] = 2704ns;

slave_timing[3][1].info_corner          = 1;
slave_timing[3][1].info_temp__j__       = 125;
slave_timing[3][1].info_i__quite_rec__  = 0.006000000;
slave_timing[3][1].info_dtr__ib__       = -1;
slave_timing[3][1].info_i__offset_rec__ = 0.000000000;
slave_timing[3][1].info_i__max_slave__  = 0.025000000;
slave_timing[3][1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][1].info_r__dsi_bus__    = 5.000;

slave_timing[3][1].t_rxd1[0][1] = 2643ns;
slave_timing[3][1].t_rxd1[1][0] = 2814ns;
slave_timing[3][1].t_rxd1[0][2] = 1993ns;
slave_timing[3][1].t_rxd1[2][0] = 3374ns;
slave_timing[3][1].t_rxd2[0][2] = 3101ns;
slave_timing[3][1].t_rxd2[2][0] = 2181ns;
slave_timing[3][1].t_rxd2[1][2] = 2435ns;
slave_timing[3][1].t_rxd2[2][1] = 2978ns;

slave_timing[3][2].info_corner          = 1;
slave_timing[3][2].info_temp__j__       = 125;
slave_timing[3][2].info_i__quite_rec__  = 0.006000000;
slave_timing[3][2].info_dtr__ib__       = 1;
slave_timing[3][2].info_i__offset_rec__ = 0.000000000;
slave_timing[3][2].info_i__max_slave__  = 0.023000000;
slave_timing[3][2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][2].info_r__dsi_bus__    = 5.000;

slave_timing[3][2].t_rxd1[0][1] = 2851ns;
slave_timing[3][2].t_rxd1[1][0] = 2638ns;
slave_timing[3][2].t_rxd1[0][2] = 2114ns;
slave_timing[3][2].t_rxd1[2][0] = 3250ns;
slave_timing[3][2].t_rxd2[0][2] = 3500ns;
slave_timing[3][2].t_rxd2[2][0] = 1878ns;
slave_timing[3][2].t_rxd2[1][2] = 3024ns;
slave_timing[3][2].t_rxd2[2][1] = 2459ns;

slave_timing[3][3].info_corner          = 1;
slave_timing[3][3].info_temp__j__       = 125;
slave_timing[3][3].info_i__quite_rec__  = 0.006000000;
slave_timing[3][3].info_dtr__ib__       = 1;
slave_timing[3][3].info_i__offset_rec__ = 0.000000000;
slave_timing[3][3].info_i__max_slave__  = 0.025000000;
slave_timing[3][3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][3].info_r__dsi_bus__    = 5.000;

slave_timing[3][3].t_rxd1[0][1] = 2737ns;
slave_timing[3][3].t_rxd1[1][0] = 2722ns;
slave_timing[3][3].t_rxd1[0][2] = 2042ns;
slave_timing[3][3].t_rxd1[2][0] = 3314ns;
slave_timing[3][3].t_rxd2[0][2] = 3263ns;
slave_timing[3][3].t_rxd2[2][0] = 2050ns;
slave_timing[3][3].t_rxd2[1][2] = 2684ns;
slave_timing[3][3].t_rxd2[2][1] = 2738ns;

slave_timing[3][4].info_corner          = 1;
slave_timing[3][4].info_temp__j__       = 125;
slave_timing[3][4].info_i__quite_rec__  = 0.006000000;
slave_timing[3][4].info_dtr__ib__       = -1;
slave_timing[3][4].info_i__offset_rec__ = 0.000000000;
slave_timing[3][4].info_i__max_slave__  = 0.023000000;
slave_timing[3][4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][4].info_r__dsi_bus__    = 5.000;

slave_timing[3][4].t_rxd1[0][1] = 2935ns;
slave_timing[3][4].t_rxd1[1][0] = 2886ns;
slave_timing[3][4].t_rxd1[0][2] = 2224ns;
slave_timing[3][4].t_rxd1[2][0] = 3470ns;
slave_timing[3][4].t_rxd2[0][2] = 3321ns;
slave_timing[3][4].t_rxd2[2][0] = 2064ns;
slave_timing[3][4].t_rxd2[1][2] = 2744ns;
slave_timing[3][4].t_rxd2[2][1] = 2730ns;

slave_timing[3][5].info_corner          = 1;
slave_timing[3][5].info_temp__j__       = 125;
slave_timing[3][5].info_i__quite_rec__  = 0.006000000;
slave_timing[3][5].info_dtr__ib__       = -1;
slave_timing[3][5].info_i__offset_rec__ = 0.000000000;
slave_timing[3][5].info_i__max_slave__  = 0.025000000;
slave_timing[3][5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][5].info_r__dsi_bus__    = 5.000;

slave_timing[3][5].t_rxd1[0][1] = 2827ns;
slave_timing[3][5].t_rxd1[1][0] = 2972ns;
slave_timing[3][5].t_rxd1[0][2] = 2160ns;
slave_timing[3][5].t_rxd1[2][0] = 3523ns;
slave_timing[3][5].t_rxd2[0][2] = 3134ns;
slave_timing[3][5].t_rxd2[2][0] = 2211ns;
slave_timing[3][5].t_rxd2[1][2] = 2497ns;
slave_timing[3][5].t_rxd2[2][1] = 2972ns;

slave_timing[3][6].info_corner          = 1;
slave_timing[3][6].info_temp__j__       = 125;
slave_timing[3][6].info_i__quite_rec__  = 0.006000000;
slave_timing[3][6].info_dtr__ib__       = 1;
slave_timing[3][6].info_i__offset_rec__ = 0.000000000;
slave_timing[3][6].info_i__max_slave__  = 0.023000000;
slave_timing[3][6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][6].info_r__dsi_bus__    = 5.000;

slave_timing[3][6].t_rxd1[0][1] = 3029ns;
slave_timing[3][6].t_rxd1[1][0] = 2795ns;
slave_timing[3][6].t_rxd1[0][2] = 2277ns;
slave_timing[3][6].t_rxd1[2][0] = 3400ns;
slave_timing[3][6].t_rxd2[0][2] = 3521ns;
slave_timing[3][6].t_rxd2[2][0] = 1911ns;
slave_timing[3][6].t_rxd2[1][2] = 3039ns;
slave_timing[3][6].t_rxd2[2][1] = 2480ns;

slave_timing[3][7].info_corner          = 1;
slave_timing[3][7].info_temp__j__       = 125;
slave_timing[3][7].info_i__quite_rec__  = 0.006000000;
slave_timing[3][7].info_dtr__ib__       = 1;
slave_timing[3][7].info_i__offset_rec__ = 0.000000000;
slave_timing[3][7].info_i__max_slave__  = 0.025000000;
slave_timing[3][7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][7].info_r__dsi_bus__    = 5.000;

slave_timing[3][7].t_rxd1[0][1] = 2915ns;
slave_timing[3][7].t_rxd1[1][0] = 2874ns;
slave_timing[3][7].t_rxd1[0][2] = 2205ns;
slave_timing[3][7].t_rxd1[2][0] = 3456ns;
slave_timing[3][7].t_rxd2[0][2] = 3287ns;
slave_timing[3][7].t_rxd2[2][0] = 2079ns;
slave_timing[3][7].t_rxd2[1][2] = 2704ns;
slave_timing[3][7].t_rxd2[2][1] = 2760ns;

slave_timing[3][8].info_corner          = 1;
slave_timing[3][8].info_temp__j__       = 125;
slave_timing[3][8].info_i__quite_rec__  = 0.003000000;
slave_timing[3][8].info_dtr__ib__       = -1;
slave_timing[3][8].info_i__offset_rec__ = 0.000000000;
slave_timing[3][8].info_i__max_slave__  = 0.023000000;
slave_timing[3][8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][8].info_r__dsi_bus__    = 5.000;

slave_timing[3][8].t_rxd1[0][1] = 2708ns;
slave_timing[3][8].t_rxd1[1][0] = 2729ns;
slave_timing[3][8].t_rxd1[0][2] = 2033ns;
slave_timing[3][8].t_rxd1[2][0] = 3317ns;
slave_timing[3][8].t_rxd2[0][2] = 3269ns;
slave_timing[3][8].t_rxd2[2][0] = 2042ns;
slave_timing[3][8].t_rxd2[1][2] = 2691ns;
slave_timing[3][8].t_rxd2[2][1] = 2684ns;

slave_timing[3][9].info_corner          = 1;
slave_timing[3][9].info_temp__j__       = 125;
slave_timing[3][9].info_i__quite_rec__  = 0.003000000;
slave_timing[3][9].info_dtr__ib__       = -1;
slave_timing[3][9].info_i__offset_rec__ = 0.000000000;
slave_timing[3][9].info_i__max_slave__  = 0.025000000;
slave_timing[3][9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][9].info_r__dsi_bus__    = 5.000;

slave_timing[3][9].t_rxd1[0][1] = 2613ns;
slave_timing[3][9].t_rxd1[1][0] = 2809ns;
slave_timing[3][9].t_rxd1[0][2] = 1966ns;
slave_timing[3][9].t_rxd1[2][0] = 3367ns;
slave_timing[3][9].t_rxd2[0][2] = 3077ns;
slave_timing[3][9].t_rxd2[2][0] = 2187ns;
slave_timing[3][9].t_rxd2[1][2] = 2411ns;
slave_timing[3][9].t_rxd2[2][1] = 3004ns;

slave_timing[3][10].info_corner          = 1;
slave_timing[3][10].info_temp__j__       = 125;
slave_timing[3][10].info_i__quite_rec__  = 0.003000000;
slave_timing[3][10].info_dtr__ib__       = 1;
slave_timing[3][10].info_i__offset_rec__ = 0.000000000;
slave_timing[3][10].info_i__max_slave__  = 0.023000000;
slave_timing[3][10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][10].info_r__dsi_bus__    = 5.000;

slave_timing[3][10].t_rxd1[0][1] = 2788ns;
slave_timing[3][10].t_rxd1[1][0] = 2641ns;
slave_timing[3][10].t_rxd1[0][2] = 2072ns;
slave_timing[3][10].t_rxd1[2][0] = 3255ns;
slave_timing[3][10].t_rxd2[0][2] = 3461ns;
slave_timing[3][10].t_rxd2[2][0] = 1884ns;
slave_timing[3][10].t_rxd2[1][2] = 2969ns;
slave_timing[3][10].t_rxd2[2][1] = 2467ns;

slave_timing[3][11].info_corner          = 1;
slave_timing[3][11].info_temp__j__       = 125;
slave_timing[3][11].info_i__quite_rec__  = 0.003000000;
slave_timing[3][11].info_dtr__ib__       = 1;
slave_timing[3][11].info_i__offset_rec__ = 0.000000000;
slave_timing[3][11].info_i__max_slave__  = 0.025000000;
slave_timing[3][11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][11].info_r__dsi_bus__    = 5.000;

slave_timing[3][11].t_rxd1[0][1] = 2676ns;
slave_timing[3][11].t_rxd1[1][0] = 2723ns;
slave_timing[3][11].t_rxd1[0][2] = 2008ns;
slave_timing[3][11].t_rxd1[2][0] = 3301ns;
slave_timing[3][11].t_rxd2[0][2] = 3231ns;
slave_timing[3][11].t_rxd2[2][0] = 2053ns;
slave_timing[3][11].t_rxd2[1][2] = 2636ns;
slave_timing[3][11].t_rxd2[2][1] = 2743ns;

slave_timing[3][12].info_corner          = 1;
slave_timing[3][12].info_temp__j__       = 125;
slave_timing[3][12].info_i__quite_rec__  = 0.003000000;
slave_timing[3][12].info_dtr__ib__       = -1;
slave_timing[3][12].info_i__offset_rec__ = 0.000000000;
slave_timing[3][12].info_i__max_slave__  = 0.023000000;
slave_timing[3][12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][12].info_r__dsi_bus__    = 5.000;

slave_timing[3][12].t_rxd1[0][1] = 2943ns;
slave_timing[3][12].t_rxd1[1][0] = 2848ns;
slave_timing[3][12].t_rxd1[0][2] = 2208ns;
slave_timing[3][12].t_rxd1[2][0] = 3466ns;
slave_timing[3][12].t_rxd2[0][2] = 3297ns;
slave_timing[3][12].t_rxd2[2][0] = 2075ns;
slave_timing[3][12].t_rxd2[1][2] = 2758ns;
slave_timing[3][12].t_rxd2[2][1] = 2707ns;

slave_timing[3][13].info_corner          = 1;
slave_timing[3][13].info_temp__j__       = 125;
slave_timing[3][13].info_i__quite_rec__  = 0.003000000;
slave_timing[3][13].info_dtr__ib__       = -1;
slave_timing[3][13].info_i__offset_rec__ = 0.000000000;
slave_timing[3][13].info_i__max_slave__  = 0.025000000;
slave_timing[3][13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][13].info_r__dsi_bus__    = 5.000;

slave_timing[3][13].t_rxd1[0][1] = 2800ns;
slave_timing[3][13].t_rxd1[1][0] = 2970ns;
slave_timing[3][13].t_rxd1[0][2] = 2137ns;
slave_timing[3][13].t_rxd1[2][0] = 3518ns;
slave_timing[3][13].t_rxd2[0][2] = 3107ns;
slave_timing[3][13].t_rxd2[2][0] = 2220ns;
slave_timing[3][13].t_rxd2[1][2] = 2438ns;
slave_timing[3][13].t_rxd2[2][1] = 3026ns;

slave_timing[3][14].info_corner          = 1;
slave_timing[3][14].info_temp__j__       = 125;
slave_timing[3][14].info_i__quite_rec__  = 0.003000000;
slave_timing[3][14].info_dtr__ib__       = 1;
slave_timing[3][14].info_i__offset_rec__ = 0.000000000;
slave_timing[3][14].info_i__max_slave__  = 0.023000000;
slave_timing[3][14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][14].info_r__dsi_bus__    = 5.000;

slave_timing[3][14].t_rxd1[0][1] = 2985ns;
slave_timing[3][14].t_rxd1[1][0] = 2794ns;
slave_timing[3][14].t_rxd1[0][2] = 2247ns;
slave_timing[3][14].t_rxd1[2][0] = 3392ns;
slave_timing[3][14].t_rxd2[0][2] = 3485ns;
slave_timing[3][14].t_rxd2[2][0] = 1910ns;
slave_timing[3][14].t_rxd2[1][2] = 2991ns;
slave_timing[3][14].t_rxd2[2][1] = 2456ns;

slave_timing[3][15].info_corner          = 1;
slave_timing[3][15].info_temp__j__       = 125;
slave_timing[3][15].info_i__quite_rec__  = 0.003000000;
slave_timing[3][15].info_dtr__ib__       = 1;
slave_timing[3][15].info_i__offset_rec__ = 0.000000000;
slave_timing[3][15].info_i__max_slave__  = 0.025000000;
slave_timing[3][15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][15].info_r__dsi_bus__    = 5.000;

slave_timing[3][15].t_rxd1[0][1] = 2871ns;
slave_timing[3][15].t_rxd1[1][0] = 2890ns;
slave_timing[3][15].t_rxd1[0][2] = 2184ns;
slave_timing[3][15].t_rxd1[2][0] = 3451ns;
slave_timing[3][15].t_rxd2[0][2] = 3257ns;
slave_timing[3][15].t_rxd2[2][0] = 2088ns;
slave_timing[3][15].t_rxd2[1][2] = 2671ns;
slave_timing[3][15].t_rxd2[2][1] = 2774ns;

slave_timing[3][16].info_corner          = 1;
slave_timing[3][16].info_temp__j__       = 125;
slave_timing[3][16].info_i__quite_rec__  = 0.000000000;
slave_timing[3][16].info_dtr__ib__       = -1;
slave_timing[3][16].info_i__offset_rec__ = 0.000000000;
slave_timing[3][16].info_i__max_slave__  = 0.023000000;
slave_timing[3][16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][16].info_r__dsi_bus__    = 5.000;

slave_timing[3][16].t_rxd1[0][1] = 2704ns;
slave_timing[3][16].t_rxd1[1][0] = 2701ns;
slave_timing[3][16].t_rxd1[0][2] = 1994ns;
slave_timing[3][16].t_rxd1[2][0] = 3289ns;
slave_timing[3][16].t_rxd2[0][2] = 3238ns;
slave_timing[3][16].t_rxd2[2][0] = 2025ns;
slave_timing[3][16].t_rxd2[1][2] = 2702ns;
slave_timing[3][16].t_rxd2[2][1] = 2686ns;

slave_timing[3][17].info_corner          = 1;
slave_timing[3][17].info_temp__j__       = 125;
slave_timing[3][17].info_i__quite_rec__  = 0.000000000;
slave_timing[3][17].info_dtr__ib__       = -1;
slave_timing[3][17].info_i__offset_rec__ = 0.000000000;
slave_timing[3][17].info_i__max_slave__  = 0.025000000;
slave_timing[3][17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][17].info_r__dsi_bus__    = 5.000;

slave_timing[3][17].t_rxd1[0][1] = 2602ns;
slave_timing[3][17].t_rxd1[1][0] = 2785ns;
slave_timing[3][17].t_rxd1[0][2] = 1956ns;
slave_timing[3][17].t_rxd1[2][0] = 3340ns;
slave_timing[3][17].t_rxd2[0][2] = 3077ns;
slave_timing[3][17].t_rxd2[2][0] = 2167ns;
slave_timing[3][17].t_rxd2[1][2] = 2416ns;
slave_timing[3][17].t_rxd2[2][1] = 2969ns;

slave_timing[3][18].info_corner          = 1;
slave_timing[3][18].info_temp__j__       = 125;
slave_timing[3][18].info_i__quite_rec__  = 0.000000000;
slave_timing[3][18].info_dtr__ib__       = 1;
slave_timing[3][18].info_i__offset_rec__ = 0.000000000;
slave_timing[3][18].info_i__max_slave__  = 0.023000000;
slave_timing[3][18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][18].info_r__dsi_bus__    = 5.000;

slave_timing[3][18].t_rxd1[0][1] = 2816ns;
slave_timing[3][18].t_rxd1[1][0] = 2585ns;
slave_timing[3][18].t_rxd1[0][2] = 2080ns;
slave_timing[3][18].t_rxd1[2][0] = 3198ns;
slave_timing[3][18].t_rxd2[0][2] = 3494ns;
slave_timing[3][18].t_rxd2[2][0] = 1823ns;
slave_timing[3][18].t_rxd2[1][2] = 3027ns;
slave_timing[3][18].t_rxd2[2][1] = 2346ns;

slave_timing[3][19].info_corner          = 1;
slave_timing[3][19].info_temp__j__       = 125;
slave_timing[3][19].info_i__quite_rec__  = 0.000000000;
slave_timing[3][19].info_dtr__ib__       = 1;
slave_timing[3][19].info_i__offset_rec__ = 0.000000000;
slave_timing[3][19].info_i__max_slave__  = 0.025000000;
slave_timing[3][19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][19].info_r__dsi_bus__    = 5.000;

slave_timing[3][19].t_rxd1[0][1] = 2703ns;
slave_timing[3][19].t_rxd1[1][0] = 2669ns;
slave_timing[3][19].t_rxd1[0][2] = 2010ns;
slave_timing[3][19].t_rxd1[2][0] = 3253ns;
slave_timing[3][19].t_rxd2[0][2] = 3251ns;
slave_timing[3][19].t_rxd2[2][0] = 2007ns;
slave_timing[3][19].t_rxd2[1][2] = 2686ns;
slave_timing[3][19].t_rxd2[2][1] = 2667ns;

slave_timing[3][20].info_corner          = 1;
slave_timing[3][20].info_temp__j__       = 125;
slave_timing[3][20].info_i__quite_rec__  = 0.000000000;
slave_timing[3][20].info_dtr__ib__       = -1;
slave_timing[3][20].info_i__offset_rec__ = 0.000000000;
slave_timing[3][20].info_i__max_slave__  = 0.023000000;
slave_timing[3][20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][20].info_r__dsi_bus__    = 5.000;

slave_timing[3][20].t_rxd1[0][1] = 2906ns;
slave_timing[3][20].t_rxd1[1][0] = 2862ns;
slave_timing[3][20].t_rxd1[0][2] = 2204ns;
slave_timing[3][20].t_rxd1[2][0] = 3434ns;
slave_timing[3][20].t_rxd2[0][2] = 3287ns;
slave_timing[3][20].t_rxd2[2][0] = 2054ns;
slave_timing[3][20].t_rxd2[1][2] = 2725ns;
slave_timing[3][20].t_rxd2[2][1] = 2714ns;

slave_timing[3][21].info_corner          = 1;
slave_timing[3][21].info_temp__j__       = 125;
slave_timing[3][21].info_i__quite_rec__  = 0.000000000;
slave_timing[3][21].info_dtr__ib__       = -1;
slave_timing[3][21].info_i__offset_rec__ = 0.000000000;
slave_timing[3][21].info_i__max_slave__  = 0.025000000;
slave_timing[3][21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][21].info_r__dsi_bus__    = 5.000;

slave_timing[3][21].t_rxd1[0][1] = 2801ns;
slave_timing[3][21].t_rxd1[1][0] = 2935ns;
slave_timing[3][21].t_rxd1[0][2] = 2146ns;
slave_timing[3][21].t_rxd1[2][0] = 3485ns;
slave_timing[3][21].t_rxd2[0][2] = 3103ns;
slave_timing[3][21].t_rxd2[2][0] = 2201ns;
slave_timing[3][21].t_rxd2[1][2] = 2443ns;
slave_timing[3][21].t_rxd2[2][1] = 2997ns;

slave_timing[3][22].info_corner          = 1;
slave_timing[3][22].info_temp__j__       = 125;
slave_timing[3][22].info_i__quite_rec__  = 0.000000000;
slave_timing[3][22].info_dtr__ib__       = 1;
slave_timing[3][22].info_i__offset_rec__ = 0.000000000;
slave_timing[3][22].info_i__max_slave__  = 0.023000000;
slave_timing[3][22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][22].info_r__dsi_bus__    = 5.000;

slave_timing[3][22].t_rxd1[0][1] = 3023ns;
slave_timing[3][22].t_rxd1[1][0] = 2737ns;
slave_timing[3][22].t_rxd1[0][2] = 2266ns;
slave_timing[3][22].t_rxd1[2][0] = 3342ns;
slave_timing[3][22].t_rxd2[0][2] = 3512ns;
slave_timing[3][22].t_rxd2[2][0] = 1850ns;
slave_timing[3][22].t_rxd2[1][2] = 3056ns;
slave_timing[3][22].t_rxd2[2][1] = 2404ns;

slave_timing[3][23].info_corner          = 1;
slave_timing[3][23].info_temp__j__       = 125;
slave_timing[3][23].info_i__quite_rec__  = 0.000000000;
slave_timing[3][23].info_dtr__ib__       = 1;
slave_timing[3][23].info_i__offset_rec__ = 0.000000000;
slave_timing[3][23].info_i__max_slave__  = 0.025000000;
slave_timing[3][23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][23].info_r__dsi_bus__    = 5.000;

slave_timing[3][23].t_rxd1[0][1] = 2908ns;
slave_timing[3][23].t_rxd1[1][0] = 2820ns;
slave_timing[3][23].t_rxd1[0][2] = 2202ns;
slave_timing[3][23].t_rxd1[2][0] = 3397ns;
slave_timing[3][23].t_rxd2[0][2] = 3274ns;
slave_timing[3][23].t_rxd2[2][0] = 2025ns;
slave_timing[3][23].t_rxd2[1][2] = 2713ns;
slave_timing[3][23].t_rxd2[2][1] = 2690ns;

slave_timing[3][24].info_corner          = 1;
slave_timing[3][24].info_temp__j__       = 125;
slave_timing[3][24].info_i__quite_rec__  = 0.040000000;
slave_timing[3][24].info_dtr__ib__       = -1;
slave_timing[3][24].info_i__offset_rec__ = 0.000000000;
slave_timing[3][24].info_i__max_slave__  = 0.023000000;
slave_timing[3][24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][24].info_r__dsi_bus__    = 5.000;

slave_timing[3][24].t_rxd1[0][1] = 2751ns;
slave_timing[3][24].t_rxd1[1][0] = 2732ns;
slave_timing[3][24].t_rxd1[0][2] = 2038ns;
slave_timing[3][24].t_rxd1[2][0] = 3344ns;
slave_timing[3][24].t_rxd2[0][2] = 3270ns;
slave_timing[3][24].t_rxd2[2][0] = 2063ns;
slave_timing[3][24].t_rxd2[1][2] = 2722ns;
slave_timing[3][24].t_rxd2[2][1] = 2705ns;

slave_timing[3][25].info_corner          = 1;
slave_timing[3][25].info_temp__j__       = 125;
slave_timing[3][25].info_i__quite_rec__  = 0.040000000;
slave_timing[3][25].info_dtr__ib__       = -1;
slave_timing[3][25].info_i__offset_rec__ = 0.000000000;
slave_timing[3][25].info_i__max_slave__  = 0.025000000;
slave_timing[3][25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][25].info_r__dsi_bus__    = 5.000;

slave_timing[3][25].t_rxd1[0][1] = 2604ns;
slave_timing[3][25].t_rxd1[1][0] = 2848ns;
slave_timing[3][25].t_rxd1[0][2] = 1968ns;
slave_timing[3][25].t_rxd1[2][0] = 3400ns;
slave_timing[3][25].t_rxd2[0][2] = 3093ns;
slave_timing[3][25].t_rxd2[2][0] = 2211ns;
slave_timing[3][25].t_rxd2[1][2] = 2401ns;
slave_timing[3][25].t_rxd2[2][1] = 3037ns;

slave_timing[3][26].info_corner          = 1;
slave_timing[3][26].info_temp__j__       = 125;
slave_timing[3][26].info_i__quite_rec__  = 0.040000000;
slave_timing[3][26].info_dtr__ib__       = 1;
slave_timing[3][26].info_i__offset_rec__ = 0.000000000;
slave_timing[3][26].info_i__max_slave__  = 0.023000000;
slave_timing[3][26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][26].info_r__dsi_bus__    = 5.000;

slave_timing[3][26].t_rxd1[0][1] = 2820ns;
slave_timing[3][26].t_rxd1[1][0] = 2665ns;
slave_timing[3][26].t_rxd1[0][2] = 2094ns;
slave_timing[3][26].t_rxd1[2][0] = 3274ns;
slave_timing[3][26].t_rxd2[0][2] = 3475ns;
slave_timing[3][26].t_rxd2[2][0] = 1902ns;
slave_timing[3][26].t_rxd2[1][2] = 2975ns;
slave_timing[3][26].t_rxd2[2][1] = 2448ns;

slave_timing[3][27].info_corner          = 1;
slave_timing[3][27].info_temp__j__       = 125;
slave_timing[3][27].info_i__quite_rec__  = 0.040000000;
slave_timing[3][27].info_dtr__ib__       = 1;
slave_timing[3][27].info_i__offset_rec__ = 0.000000000;
slave_timing[3][27].info_i__max_slave__  = 0.025000000;
slave_timing[3][27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][27].info_r__dsi_bus__    = 5.000;

slave_timing[3][27].t_rxd1[0][1] = 2707ns;
slave_timing[3][27].t_rxd1[1][0] = 2746ns;
slave_timing[3][27].t_rxd1[0][2] = 2023ns;
slave_timing[3][27].t_rxd1[2][0] = 3327ns;
slave_timing[3][27].t_rxd2[0][2] = 3248ns;
slave_timing[3][27].t_rxd2[2][0] = 2071ns;
slave_timing[3][27].t_rxd2[1][2] = 2689ns;
slave_timing[3][27].t_rxd2[2][1] = 2736ns;

slave_timing[3][28].info_corner          = 1;
slave_timing[3][28].info_temp__j__       = 125;
slave_timing[3][28].info_i__quite_rec__  = 0.040000000;
slave_timing[3][28].info_dtr__ib__       = -1;
slave_timing[3][28].info_i__offset_rec__ = 0.000000000;
slave_timing[3][28].info_i__max_slave__  = 0.023000000;
slave_timing[3][28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][28].info_r__dsi_bus__    = 5.000;

slave_timing[3][28].t_rxd1[0][1] = 2808ns;
slave_timing[3][28].t_rxd1[1][0] = 2868ns;
slave_timing[3][28].t_rxd1[0][2] = 2126ns;
slave_timing[3][28].t_rxd1[2][0] = 3441ns;
slave_timing[3][28].t_rxd2[0][2] = 3303ns;
slave_timing[3][28].t_rxd2[2][0] = 2095ns;
slave_timing[3][28].t_rxd2[1][2] = 2723ns;
slave_timing[3][28].t_rxd2[2][1] = 2777ns;

slave_timing[3][29].info_corner          = 1;
slave_timing[3][29].info_temp__j__       = 125;
slave_timing[3][29].info_i__quite_rec__  = 0.040000000;
slave_timing[3][29].info_dtr__ib__       = -1;
slave_timing[3][29].info_i__offset_rec__ = 0.000000000;
slave_timing[3][29].info_i__max_slave__  = 0.025000000;
slave_timing[3][29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][29].info_r__dsi_bus__    = 5.000;

slave_timing[3][29].t_rxd1[0][1] = 2747ns;
slave_timing[3][29].t_rxd1[1][0] = 2912ns;
slave_timing[3][29].t_rxd1[0][2] = 2089ns;
slave_timing[3][29].t_rxd1[2][0] = 3463ns;
slave_timing[3][29].t_rxd2[0][2] = 3143ns;
slave_timing[3][29].t_rxd2[2][0] = 2215ns;
slave_timing[3][29].t_rxd2[1][2] = 2479ns;
slave_timing[3][29].t_rxd2[2][1] = 3018ns;

slave_timing[3][30].info_corner          = 1;
slave_timing[3][30].info_temp__j__       = 125;
slave_timing[3][30].info_i__quite_rec__  = 0.040000000;
slave_timing[3][30].info_dtr__ib__       = 1;
slave_timing[3][30].info_i__offset_rec__ = 0.000000000;
slave_timing[3][30].info_i__max_slave__  = 0.023000000;
slave_timing[3][30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][30].info_r__dsi_bus__    = 5.000;

slave_timing[3][30].t_rxd1[0][1] = 2922ns;
slave_timing[3][30].t_rxd1[1][0] = 2757ns;
slave_timing[3][30].t_rxd1[0][2] = 2185ns;
slave_timing[3][30].t_rxd1[2][0] = 3361ns;
slave_timing[3][30].t_rxd2[0][2] = 3509ns;
slave_timing[3][30].t_rxd2[2][0] = 1935ns;
slave_timing[3][30].t_rxd2[1][2] = 3008ns;
slave_timing[3][30].t_rxd2[2][1] = 2525ns;

slave_timing[3][31].info_corner          = 1;
slave_timing[3][31].info_temp__j__       = 125;
slave_timing[3][31].info_i__quite_rec__  = 0.040000000;
slave_timing[3][31].info_dtr__ib__       = 1;
slave_timing[3][31].info_i__offset_rec__ = 0.000000000;
slave_timing[3][31].info_i__max_slave__  = 0.025000000;
slave_timing[3][31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][31].info_r__dsi_bus__    = 5.000;

slave_timing[3][31].t_rxd1[0][1] = 2809ns;
slave_timing[3][31].t_rxd1[1][0] = 2844ns;
slave_timing[3][31].t_rxd1[0][2] = 2122ns;
slave_timing[3][31].t_rxd1[2][0] = 3419ns;
slave_timing[3][31].t_rxd2[0][2] = 3285ns;
slave_timing[3][31].t_rxd2[2][0] = 2108ns;
slave_timing[3][31].t_rxd2[1][2] = 2687ns;
slave_timing[3][31].t_rxd2[2][1] = 2801ns;

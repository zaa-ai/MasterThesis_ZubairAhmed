`define SVN_REVISION 16'd1178


slave_timing[0][64+0].info_corner          = 3;
slave_timing[0][64+0].info_temp__j__       = 125;
slave_timing[0][64+0].info_i__quite_rec__  = 0.006000000;
slave_timing[0][64+0].info_dtr__ib__       = -1;
slave_timing[0][64+0].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+0].info_i__max_slave__  = 0.023000000;
slave_timing[0][64+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][64+0].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+0].t_rxd1[0][1] = 1091ns;
slave_timing[0][64+0].t_rxd1[1][0] = 1092ns;
slave_timing[0][64+0].t_rxd1[0][2] = 804ns;
slave_timing[0][64+0].t_rxd1[2][0] = 1351ns;
slave_timing[0][64+0].t_rxd2[0][2] = 1322ns;
slave_timing[0][64+0].t_rxd2[2][0] = 818ns;
slave_timing[0][64+0].t_rxd2[1][2] = 1086ns;
slave_timing[0][64+0].t_rxd2[2][1] = 1088ns;

slave_timing[0][64+1].info_corner          = 3;
slave_timing[0][64+1].info_temp__j__       = 125;
slave_timing[0][64+1].info_i__quite_rec__  = 0.006000000;
slave_timing[0][64+1].info_dtr__ib__       = -1;
slave_timing[0][64+1].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+1].info_i__max_slave__  = 0.025000000;
slave_timing[0][64+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][64+1].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+1].t_rxd1[0][1] = 1046ns;
slave_timing[0][64+1].t_rxd1[1][0] = 1124ns;
slave_timing[0][64+1].t_rxd1[0][2] = 787ns;
slave_timing[0][64+1].t_rxd1[2][0] = 1380ns;
slave_timing[0][64+1].t_rxd2[0][2] = 1241ns;
slave_timing[0][64+1].t_rxd2[2][0] = 871ns;
slave_timing[0][64+1].t_rxd2[1][2] = 962ns;
slave_timing[0][64+1].t_rxd2[2][1] = 1214ns;

slave_timing[0][64+2].info_corner          = 3;
slave_timing[0][64+2].info_temp__j__       = 125;
slave_timing[0][64+2].info_i__quite_rec__  = 0.006000000;
slave_timing[0][64+2].info_dtr__ib__       = 1;
slave_timing[0][64+2].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+2].info_i__max_slave__  = 0.023000000;
slave_timing[0][64+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][64+2].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+2].t_rxd1[0][1] = 1102ns;
slave_timing[0][64+2].t_rxd1[1][0] = 1047ns;
slave_timing[0][64+2].t_rxd1[0][2] = 812ns;
slave_timing[0][64+2].t_rxd1[2][0] = 1305ns;
slave_timing[0][64+2].t_rxd2[0][2] = 1405ns;
slave_timing[0][64+2].t_rxd2[2][0] = 768ns;
slave_timing[0][64+2].t_rxd2[1][2] = 1181ns;
slave_timing[0][64+2].t_rxd2[2][1] = 989ns;

slave_timing[0][64+3].info_corner          = 3;
slave_timing[0][64+3].info_temp__j__       = 125;
slave_timing[0][64+3].info_i__quite_rec__  = 0.006000000;
slave_timing[0][64+3].info_dtr__ib__       = 1;
slave_timing[0][64+3].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+3].info_i__max_slave__  = 0.025000000;
slave_timing[0][64+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][64+3].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+3].t_rxd1[0][1] = 1053ns;
slave_timing[0][64+3].t_rxd1[1][0] = 1080ns;
slave_timing[0][64+3].t_rxd1[0][2] = 789ns;
slave_timing[0][64+3].t_rxd1[2][0] = 1330ns;
slave_timing[0][64+3].t_rxd2[0][2] = 1286ns;
slave_timing[0][64+3].t_rxd2[2][0] = 824ns;
slave_timing[0][64+3].t_rxd2[1][2] = 1040ns;
slave_timing[0][64+3].t_rxd2[2][1] = 1105ns;

slave_timing[0][64+4].info_corner          = 3;
slave_timing[0][64+4].info_temp__j__       = 125;
slave_timing[0][64+4].info_i__quite_rec__  = 0.006000000;
slave_timing[0][64+4].info_dtr__ib__       = -1;
slave_timing[0][64+4].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+4].info_i__max_slave__  = 0.023000000;
slave_timing[0][64+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][64+4].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+4].t_rxd1[0][1] = 1294ns;
slave_timing[0][64+4].t_rxd1[1][0] = 1239ns;
slave_timing[0][64+4].t_rxd1[0][2] = 953ns;
slave_timing[0][64+4].t_rxd1[2][0] = 1489ns;
slave_timing[0][64+4].t_rxd2[0][2] = 1410ns;
slave_timing[0][64+4].t_rxd2[2][0] = 858ns;
slave_timing[0][64+4].t_rxd2[1][2] = 1115ns;
slave_timing[0][64+4].t_rxd2[2][1] = 1119ns;

slave_timing[0][64+5].info_corner          = 3;
slave_timing[0][64+5].info_temp__j__       = 125;
slave_timing[0][64+5].info_i__quite_rec__  = 0.006000000;
slave_timing[0][64+5].info_dtr__ib__       = -1;
slave_timing[0][64+5].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+5].info_i__max_slave__  = 0.025000000;
slave_timing[0][64+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][64+5].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+5].t_rxd1[0][1] = 1237ns;
slave_timing[0][64+5].t_rxd1[1][0] = 1272ns;
slave_timing[0][64+5].t_rxd1[0][2] = 926ns;
slave_timing[0][64+5].t_rxd1[2][0] = 1515ns;
slave_timing[0][64+5].t_rxd2[0][2] = 1313ns;
slave_timing[0][64+5].t_rxd2[2][0] = 910ns;
slave_timing[0][64+5].t_rxd2[1][2] = 997ns;
slave_timing[0][64+5].t_rxd2[2][1] = 1235ns;

slave_timing[0][64+6].info_corner          = 3;
slave_timing[0][64+6].info_temp__j__       = 125;
slave_timing[0][64+6].info_i__quite_rec__  = 0.006000000;
slave_timing[0][64+6].info_dtr__ib__       = 1;
slave_timing[0][64+6].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+6].info_i__max_slave__  = 0.023000000;
slave_timing[0][64+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][64+6].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+6].t_rxd1[0][1] = 1298ns;
slave_timing[0][64+6].t_rxd1[1][0] = 1184ns;
slave_timing[0][64+6].t_rxd1[0][2] = 948ns;
slave_timing[0][64+6].t_rxd1[2][0] = 1429ns;
slave_timing[0][64+6].t_rxd2[0][2] = 1469ns;
slave_timing[0][64+6].t_rxd2[2][0] = 801ns;
slave_timing[0][64+6].t_rxd2[1][2] = 1203ns;
slave_timing[0][64+6].t_rxd2[2][1] = 1019ns;

slave_timing[0][64+7].info_corner          = 3;
slave_timing[0][64+7].info_temp__j__       = 125;
slave_timing[0][64+7].info_i__quite_rec__  = 0.006000000;
slave_timing[0][64+7].info_dtr__ib__       = 1;
slave_timing[0][64+7].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+7].info_i__max_slave__  = 0.025000000;
slave_timing[0][64+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][64+7].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+7].t_rxd1[0][1] = 1240ns;
slave_timing[0][64+7].t_rxd1[1][0] = 1216ns;
slave_timing[0][64+7].t_rxd1[0][2] = 920ns;
slave_timing[0][64+7].t_rxd1[2][0] = 1458ns;
slave_timing[0][64+7].t_rxd2[0][2] = 1350ns;
slave_timing[0][64+7].t_rxd2[2][0] = 860ns;
slave_timing[0][64+7].t_rxd2[1][2] = 1067ns;
slave_timing[0][64+7].t_rxd2[2][1] = 1131ns;

slave_timing[0][64+8].info_corner          = 3;
slave_timing[0][64+8].info_temp__j__       = 125;
slave_timing[0][64+8].info_i__quite_rec__  = 0.003000000;
slave_timing[0][64+8].info_dtr__ib__       = -1;
slave_timing[0][64+8].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+8].info_i__max_slave__  = 0.023000000;
slave_timing[0][64+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][64+8].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+8].t_rxd1[0][1] = 1047ns;
slave_timing[0][64+8].t_rxd1[1][0] = 1073ns;
slave_timing[0][64+8].t_rxd1[0][2] = 786ns;
slave_timing[0][64+8].t_rxd1[2][0] = 1315ns;
slave_timing[0][64+8].t_rxd2[0][2] = 1288ns;
slave_timing[0][64+8].t_rxd2[2][0] = 805ns;
slave_timing[0][64+8].t_rxd2[1][2] = 1054ns;
slave_timing[0][64+8].t_rxd2[2][1] = 1071ns;

slave_timing[0][64+9].info_corner          = 3;
slave_timing[0][64+9].info_temp__j__       = 125;
slave_timing[0][64+9].info_i__quite_rec__  = 0.003000000;
slave_timing[0][64+9].info_dtr__ib__       = -1;
slave_timing[0][64+9].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+9].info_i__max_slave__  = 0.025000000;
slave_timing[0][64+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][64+9].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+9].t_rxd1[0][1] = 1004ns;
slave_timing[0][64+9].t_rxd1[1][0] = 1104ns;
slave_timing[0][64+9].t_rxd1[0][2] = 762ns;
slave_timing[0][64+9].t_rxd1[2][0] = 1342ns;
slave_timing[0][64+9].t_rxd2[0][2] = 1197ns;
slave_timing[0][64+9].t_rxd2[2][0] = 857ns;
slave_timing[0][64+9].t_rxd2[1][2] = 935ns;
slave_timing[0][64+9].t_rxd2[2][1] = 1189ns;

slave_timing[0][64+10].info_corner          = 3;
slave_timing[0][64+10].info_temp__j__       = 125;
slave_timing[0][64+10].info_i__quite_rec__  = 0.003000000;
slave_timing[0][64+10].info_dtr__ib__       = 1;
slave_timing[0][64+10].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+10].info_i__max_slave__  = 0.023000000;
slave_timing[0][64+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][64+10].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+10].t_rxd1[0][1] = 1072ns;
slave_timing[0][64+10].t_rxd1[1][0] = 1013ns;
slave_timing[0][64+10].t_rxd1[0][2] = 791ns;
slave_timing[0][64+10].t_rxd1[2][0] = 1249ns;
slave_timing[0][64+10].t_rxd2[0][2] = 1365ns;
slave_timing[0][64+10].t_rxd2[2][0] = 744ns;
slave_timing[0][64+10].t_rxd2[1][2] = 1160ns;
slave_timing[0][64+10].t_rxd2[2][1] = 959ns;

slave_timing[0][64+11].info_corner          = 3;
slave_timing[0][64+11].info_temp__j__       = 125;
slave_timing[0][64+11].info_i__quite_rec__  = 0.003000000;
slave_timing[0][64+11].info_dtr__ib__       = 1;
slave_timing[0][64+11].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+11].info_i__max_slave__  = 0.025000000;
slave_timing[0][64+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][64+11].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+11].t_rxd1[0][1] = 1025ns;
slave_timing[0][64+11].t_rxd1[1][0] = 1042ns;
slave_timing[0][64+11].t_rxd1[0][2] = 770ns;
slave_timing[0][64+11].t_rxd1[2][0] = 1279ns;
slave_timing[0][64+11].t_rxd2[0][2] = 1250ns;
slave_timing[0][64+11].t_rxd2[2][0] = 805ns;
slave_timing[0][64+11].t_rxd2[1][2] = 1023ns;
slave_timing[0][64+11].t_rxd2[2][1] = 1069ns;

slave_timing[0][64+12].info_corner          = 3;
slave_timing[0][64+12].info_temp__j__       = 125;
slave_timing[0][64+12].info_i__quite_rec__  = 0.003000000;
slave_timing[0][64+12].info_dtr__ib__       = -1;
slave_timing[0][64+12].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+12].info_i__max_slave__  = 0.023000000;
slave_timing[0][64+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][64+12].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+12].t_rxd1[0][1] = 1267ns;
slave_timing[0][64+12].t_rxd1[1][0] = 1220ns;
slave_timing[0][64+12].t_rxd1[0][2] = 937ns;
slave_timing[0][64+12].t_rxd1[2][0] = 1452ns;
slave_timing[0][64+12].t_rxd2[0][2] = 1358ns;
slave_timing[0][64+12].t_rxd2[2][0] = 846ns;
slave_timing[0][64+12].t_rxd2[1][2] = 1100ns;
slave_timing[0][64+12].t_rxd2[2][1] = 1085ns;

slave_timing[0][64+13].info_corner          = 3;
slave_timing[0][64+13].info_temp__j__       = 125;
slave_timing[0][64+13].info_i__quite_rec__  = 0.003000000;
slave_timing[0][64+13].info_dtr__ib__       = -1;
slave_timing[0][64+13].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+13].info_i__max_slave__  = 0.025000000;
slave_timing[0][64+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][64+13].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+13].t_rxd1[0][1] = 1213ns;
slave_timing[0][64+13].t_rxd1[1][0] = 1247ns;
slave_timing[0][64+13].t_rxd1[0][2] = 910ns;
slave_timing[0][64+13].t_rxd1[2][0] = 1475ns;
slave_timing[0][64+13].t_rxd2[0][2] = 1270ns;
slave_timing[0][64+13].t_rxd2[2][0] = 893ns;
slave_timing[0][64+13].t_rxd2[1][2] = 970ns;
slave_timing[0][64+13].t_rxd2[2][1] = 1197ns;

slave_timing[0][64+14].info_corner          = 3;
slave_timing[0][64+14].info_temp__j__       = 125;
slave_timing[0][64+14].info_i__quite_rec__  = 0.003000000;
slave_timing[0][64+14].info_dtr__ib__       = 1;
slave_timing[0][64+14].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+14].info_i__max_slave__  = 0.023000000;
slave_timing[0][64+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][64+14].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+14].t_rxd1[0][1] = 1290ns;
slave_timing[0][64+14].t_rxd1[1][0] = 1144ns;
slave_timing[0][64+14].t_rxd1[0][2] = 943ns;
slave_timing[0][64+14].t_rxd1[2][0] = 1377ns;
slave_timing[0][64+14].t_rxd2[0][2] = 1428ns;
slave_timing[0][64+14].t_rxd2[2][0] = 782ns;
slave_timing[0][64+14].t_rxd2[1][2] = 1181ns;
slave_timing[0][64+14].t_rxd2[2][1] = 990ns;

slave_timing[0][64+15].info_corner          = 3;
slave_timing[0][64+15].info_temp__j__       = 125;
slave_timing[0][64+15].info_i__quite_rec__  = 0.003000000;
slave_timing[0][64+15].info_dtr__ib__       = 1;
slave_timing[0][64+15].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+15].info_i__max_slave__  = 0.025000000;
slave_timing[0][64+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][64+15].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+15].t_rxd1[0][1] = 1233ns;
slave_timing[0][64+15].t_rxd1[1][0] = 1178ns;
slave_timing[0][64+15].t_rxd1[0][2] = 915ns;
slave_timing[0][64+15].t_rxd1[2][0] = 1401ns;
slave_timing[0][64+15].t_rxd2[0][2] = 1314ns;
slave_timing[0][64+15].t_rxd2[2][0] = 839ns;
slave_timing[0][64+15].t_rxd2[1][2] = 1050ns;
slave_timing[0][64+15].t_rxd2[2][1] = 1095ns;

slave_timing[0][64+16].info_corner          = 3;
slave_timing[0][64+16].info_temp__j__       = 125;
slave_timing[0][64+16].info_i__quite_rec__  = 0.000000000;
slave_timing[0][64+16].info_dtr__ib__       = -1;
slave_timing[0][64+16].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+16].info_i__max_slave__  = 0.023000000;
slave_timing[0][64+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][64+16].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+16].t_rxd1[0][1] = 1027ns;
slave_timing[0][64+16].t_rxd1[1][0] = 1035ns;
slave_timing[0][64+16].t_rxd1[0][2] = 771ns;
slave_timing[0][64+16].t_rxd1[2][0] = 1257ns;
slave_timing[0][64+16].t_rxd2[0][2] = 1247ns;
slave_timing[0][64+16].t_rxd2[2][0] = 787ns;
slave_timing[0][64+16].t_rxd2[1][2] = 1032ns;
slave_timing[0][64+16].t_rxd2[2][1] = 1038ns;

slave_timing[0][64+17].info_corner          = 3;
slave_timing[0][64+17].info_temp__j__       = 125;
slave_timing[0][64+17].info_i__quite_rec__  = 0.000000000;
slave_timing[0][64+17].info_dtr__ib__       = -1;
slave_timing[0][64+17].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+17].info_i__max_slave__  = 0.025000000;
slave_timing[0][64+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][64+17].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+17].t_rxd1[0][1] = 986ns;
slave_timing[0][64+17].t_rxd1[1][0] = 1063ns;
slave_timing[0][64+17].t_rxd1[0][2] = 748ns;
slave_timing[0][64+17].t_rxd1[2][0] = 1278ns;
slave_timing[0][64+17].t_rxd2[0][2] = 1162ns;
slave_timing[0][64+17].t_rxd2[2][0] = 833ns;
slave_timing[0][64+17].t_rxd2[1][2] = 921ns;
slave_timing[0][64+17].t_rxd2[2][1] = 1152ns;

slave_timing[0][64+18].info_corner          = 3;
slave_timing[0][64+18].info_temp__j__       = 125;
slave_timing[0][64+18].info_i__quite_rec__  = 0.000000000;
slave_timing[0][64+18].info_dtr__ib__       = 1;
slave_timing[0][64+18].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+18].info_i__max_slave__  = 0.023000000;
slave_timing[0][64+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][64+18].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+18].t_rxd1[0][1] = 1054ns;
slave_timing[0][64+18].t_rxd1[1][0] = 977ns;
slave_timing[0][64+18].t_rxd1[0][2] = 779ns;
slave_timing[0][64+18].t_rxd1[2][0] = 1200ns;
slave_timing[0][64+18].t_rxd2[0][2] = 1317ns;
slave_timing[0][64+18].t_rxd2[2][0] = 727ns;
slave_timing[0][64+18].t_rxd2[1][2] = 1125ns;
slave_timing[0][64+18].t_rxd2[2][1] = 930ns;

slave_timing[0][64+19].info_corner          = 3;
slave_timing[0][64+19].info_temp__j__       = 125;
slave_timing[0][64+19].info_i__quite_rec__  = 0.000000000;
slave_timing[0][64+19].info_dtr__ib__       = 1;
slave_timing[0][64+19].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+19].info_i__max_slave__  = 0.025000000;
slave_timing[0][64+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][64+19].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+19].t_rxd1[0][1] = 1007ns;
slave_timing[0][64+19].t_rxd1[1][0] = 1009ns;
slave_timing[0][64+19].t_rxd1[0][2] = 757ns;
slave_timing[0][64+19].t_rxd1[2][0] = 1223ns;
slave_timing[0][64+19].t_rxd2[0][2] = 1208ns;
slave_timing[0][64+19].t_rxd2[2][0] = 780ns;
slave_timing[0][64+19].t_rxd2[1][2] = 997ns;
slave_timing[0][64+19].t_rxd2[2][1] = 1032ns;

slave_timing[0][64+20].info_corner          = 3;
slave_timing[0][64+20].info_temp__j__       = 125;
slave_timing[0][64+20].info_i__quite_rec__  = 0.000000000;
slave_timing[0][64+20].info_dtr__ib__       = -1;
slave_timing[0][64+20].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+20].info_i__max_slave__  = 0.023000000;
slave_timing[0][64+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][64+20].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+20].t_rxd1[0][1] = 1269ns;
slave_timing[0][64+20].t_rxd1[1][0] = 1174ns;
slave_timing[0][64+20].t_rxd1[0][2] = 933ns;
slave_timing[0][64+20].t_rxd1[2][0] = 1381ns;
slave_timing[0][64+20].t_rxd2[0][2] = 1313ns;
slave_timing[0][64+20].t_rxd2[2][0] = 823ns;
slave_timing[0][64+20].t_rxd2[1][2] = 1051ns;
slave_timing[0][64+20].t_rxd2[2][1] = 1064ns;

slave_timing[0][64+21].info_corner          = 3;
slave_timing[0][64+21].info_temp__j__       = 125;
slave_timing[0][64+21].info_i__quite_rec__  = 0.000000000;
slave_timing[0][64+21].info_dtr__ib__       = -1;
slave_timing[0][64+21].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+21].info_i__max_slave__  = 0.025000000;
slave_timing[0][64+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][64+21].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+21].t_rxd1[0][1] = 1212ns;
slave_timing[0][64+21].t_rxd1[1][0] = 1201ns;
slave_timing[0][64+21].t_rxd1[0][2] = 908ns;
slave_timing[0][64+21].t_rxd1[2][0] = 1404ns;
slave_timing[0][64+21].t_rxd2[0][2] = 1233ns;
slave_timing[0][64+21].t_rxd2[2][0] = 871ns;
slave_timing[0][64+21].t_rxd2[1][2] = 946ns;
slave_timing[0][64+21].t_rxd2[2][1] = 1170ns;

slave_timing[0][64+22].info_corner          = 3;
slave_timing[0][64+22].info_temp__j__       = 125;
slave_timing[0][64+22].info_i__quite_rec__  = 0.000000000;
slave_timing[0][64+22].info_dtr__ib__       = 1;
slave_timing[0][64+22].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+22].info_i__max_slave__  = 0.023000000;
slave_timing[0][64+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][64+22].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+22].t_rxd1[0][1] = 1298ns;
slave_timing[0][64+22].t_rxd1[1][0] = 1109ns;
slave_timing[0][64+22].t_rxd1[0][2] = 943ns;
slave_timing[0][64+22].t_rxd1[2][0] = 1317ns;
slave_timing[0][64+22].t_rxd2[0][2] = 1376ns;
slave_timing[0][64+22].t_rxd2[2][0] = 758ns;
slave_timing[0][64+22].t_rxd2[1][2] = 1146ns;
slave_timing[0][64+22].t_rxd2[2][1] = 956ns;

slave_timing[0][64+23].info_corner          = 3;
slave_timing[0][64+23].info_temp__j__       = 125;
slave_timing[0][64+23].info_i__quite_rec__  = 0.000000000;
slave_timing[0][64+23].info_dtr__ib__       = 1;
slave_timing[0][64+23].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+23].info_i__max_slave__  = 0.025000000;
slave_timing[0][64+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][64+23].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+23].t_rxd1[0][1] = 1238ns;
slave_timing[0][64+23].t_rxd1[1][0] = 1138ns;
slave_timing[0][64+23].t_rxd1[0][2] = 915ns;
slave_timing[0][64+23].t_rxd1[2][0] = 1340ns;
slave_timing[0][64+23].t_rxd2[0][2] = 1272ns;
slave_timing[0][64+23].t_rxd2[2][0] = 814ns;
slave_timing[0][64+23].t_rxd2[1][2] = 1023ns;
slave_timing[0][64+23].t_rxd2[2][1] = 1058ns;

slave_timing[0][64+24].info_corner          = 3;
slave_timing[0][64+24].info_temp__j__       = 125;
slave_timing[0][64+24].info_i__quite_rec__  = 0.040000000;
slave_timing[0][64+24].info_dtr__ib__       = -1;
slave_timing[0][64+24].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+24].info_i__max_slave__  = 0.023000000;
slave_timing[0][64+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][64+24].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+24].t_rxd1[0][1] = 1113ns;
slave_timing[0][64+24].t_rxd1[1][0] = 1126ns;
slave_timing[0][64+24].t_rxd1[0][2] = 829ns;
slave_timing[0][64+24].t_rxd1[2][0] = 1384ns;
slave_timing[0][64+24].t_rxd2[0][2] = 1400ns;
slave_timing[0][64+24].t_rxd2[2][0] = 863ns;
slave_timing[0][64+24].t_rxd2[1][2] = 1117ns;
slave_timing[0][64+24].t_rxd2[2][1] = 1120ns;

slave_timing[0][64+25].info_corner          = 3;
slave_timing[0][64+25].info_temp__j__       = 125;
slave_timing[0][64+25].info_i__quite_rec__  = 0.040000000;
slave_timing[0][64+25].info_dtr__ib__       = -1;
slave_timing[0][64+25].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+25].info_i__max_slave__  = 0.025000000;
slave_timing[0][64+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][64+25].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+25].t_rxd1[0][1] = 1066ns;
slave_timing[0][64+25].t_rxd1[1][0] = 1158ns;
slave_timing[0][64+25].t_rxd1[0][2] = 806ns;
slave_timing[0][64+25].t_rxd1[2][0] = 1415ns;
slave_timing[0][64+25].t_rxd2[0][2] = 1313ns;
slave_timing[0][64+25].t_rxd2[2][0] = 916ns;
slave_timing[0][64+25].t_rxd2[1][2] = 1003ns;
slave_timing[0][64+25].t_rxd2[2][1] = 1253ns;

slave_timing[0][64+26].info_corner          = 3;
slave_timing[0][64+26].info_temp__j__       = 125;
slave_timing[0][64+26].info_i__quite_rec__  = 0.040000000;
slave_timing[0][64+26].info_dtr__ib__       = 1;
slave_timing[0][64+26].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+26].info_i__max_slave__  = 0.023000000;
slave_timing[0][64+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][64+26].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+26].t_rxd1[0][1] = 1145ns;
slave_timing[0][64+26].t_rxd1[1][0] = 1099ns;
slave_timing[0][64+26].t_rxd1[0][2] = 841ns;
slave_timing[0][64+26].t_rxd1[2][0] = 1361ns;
slave_timing[0][64+26].t_rxd2[0][2] = 1488ns;
slave_timing[0][64+26].t_rxd2[2][0] = 818ns;
slave_timing[0][64+26].t_rxd2[1][2] = 1224ns;
slave_timing[0][64+26].t_rxd2[2][1] = 1036ns;

slave_timing[0][64+27].info_corner          = 3;
slave_timing[0][64+27].info_temp__j__       = 125;
slave_timing[0][64+27].info_i__quite_rec__  = 0.040000000;
slave_timing[0][64+27].info_dtr__ib__       = 1;
slave_timing[0][64+27].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+27].info_i__max_slave__  = 0.025000000;
slave_timing[0][64+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][64+27].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+27].t_rxd1[0][1] = 1093ns;
slave_timing[0][64+27].t_rxd1[1][0] = 1133ns;
slave_timing[0][64+27].t_rxd1[0][2] = 820ns;
slave_timing[0][64+27].t_rxd1[2][0] = 1395ns;
slave_timing[0][64+27].t_rxd2[0][2] = 1381ns;
slave_timing[0][64+27].t_rxd2[2][0] = 879ns;
slave_timing[0][64+27].t_rxd2[1][2] = 1095ns;
slave_timing[0][64+27].t_rxd2[2][1] = 1163ns;

slave_timing[0][64+28].info_corner          = 3;
slave_timing[0][64+28].info_temp__j__       = 125;
slave_timing[0][64+28].info_i__quite_rec__  = 0.040000000;
slave_timing[0][64+28].info_dtr__ib__       = -1;
slave_timing[0][64+28].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+28].info_i__max_slave__  = 0.023000000;
slave_timing[0][64+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][64+28].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+28].t_rxd1[0][1] = 1215ns;
slave_timing[0][64+28].t_rxd1[1][0] = 1209ns;
slave_timing[0][64+28].t_rxd1[0][2] = 923ns;
slave_timing[0][64+28].t_rxd1[2][0] = 1442ns;
slave_timing[0][64+28].t_rxd2[0][2] = 1509ns;
slave_timing[0][64+28].t_rxd2[2][0] = 1133ns;
slave_timing[0][64+28].t_rxd2[1][2] = 1208ns;
slave_timing[0][64+28].t_rxd2[2][1] = 1488ns;

slave_timing[0][64+29].info_corner          = 3;
slave_timing[0][64+29].info_temp__j__       = 125;
slave_timing[0][64+29].info_i__quite_rec__  = 0.040000000;
slave_timing[0][64+29].info_dtr__ib__       = -1;
slave_timing[0][64+29].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+29].info_i__max_slave__  = 0.025000000;
slave_timing[0][64+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][64+29].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+29].t_rxd1[0][1] = 1169ns;
slave_timing[0][64+29].t_rxd1[1][0] = 1241ns;
slave_timing[0][64+29].t_rxd1[0][2] = 898ns;
slave_timing[0][64+29].t_rxd1[2][0] = 1528ns;
slave_timing[0][64+29].t_rxd2[0][2] = 1440ns;
slave_timing[0][64+29].t_rxd2[2][0] = 1230ns;
slave_timing[0][64+29].t_rxd2[1][2] = 1098ns;
slave_timing[0][64+29].t_rxd2[2][1] = 1725ns;

slave_timing[0][64+30].info_corner          = 3;
slave_timing[0][64+30].info_temp__j__       = 125;
slave_timing[0][64+30].info_i__quite_rec__  = 0.040000000;
slave_timing[0][64+30].info_dtr__ib__       = 1;
slave_timing[0][64+30].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+30].info_i__max_slave__  = 0.023000000;
slave_timing[0][64+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][64+30].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+30].t_rxd1[0][1] = 1242ns;
slave_timing[0][64+30].t_rxd1[1][0] = 1176ns;
slave_timing[0][64+30].t_rxd1[0][2] = 935ns;
slave_timing[0][64+30].t_rxd1[2][0] = 1399ns;
slave_timing[0][64+30].t_rxd2[0][2] = 1600ns;
slave_timing[0][64+30].t_rxd2[2][0] = 1065ns;
slave_timing[0][64+30].t_rxd2[1][2] = 1320ns;
slave_timing[0][64+30].t_rxd2[2][1] = 1365ns;

slave_timing[0][64+31].info_corner          = 3;
slave_timing[0][64+31].info_temp__j__       = 125;
slave_timing[0][64+31].info_i__quite_rec__  = 0.040000000;
slave_timing[0][64+31].info_dtr__ib__       = 1;
slave_timing[0][64+31].info_i__offset_rec__ = 0.000000000;
slave_timing[0][64+31].info_i__max_slave__  = 0.025000000;
slave_timing[0][64+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][64+31].info_r__dsi_bus__    = 5.000;

slave_timing[0][64+31].t_rxd1[0][1] = 1192ns;
slave_timing[0][64+31].t_rxd1[1][0] = 1212ns;
slave_timing[0][64+31].t_rxd1[0][2] = 909ns;
slave_timing[0][64+31].t_rxd1[2][0] = 1481ns;
slave_timing[0][64+31].t_rxd2[0][2] = 1510ns;
slave_timing[0][64+31].t_rxd2[2][0] = 1165ns;
slave_timing[0][64+31].t_rxd2[1][2] = 1199ns;
slave_timing[0][64+31].t_rxd2[2][1] = 1584ns;


slave_timing[2][96+0].info_corner          = 4;
slave_timing[2][96+0].info_temp__j__       = 125;
slave_timing[2][96+0].info_i__quite_rec__  = 0.006000000;
slave_timing[2][96+0].info_dtr__ib__       = -1;
slave_timing[2][96+0].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+0].info_i__max_slave__  = 0.023000000;
slave_timing[2][96+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][96+0].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+0].t_rxd1[0][1] = 2194ns;
slave_timing[2][96+0].t_rxd1[1][0] = 2156ns;
slave_timing[2][96+0].t_rxd1[0][2] = 1655ns;
slave_timing[2][96+0].t_rxd1[2][0] = 2640ns;
slave_timing[2][96+0].t_rxd2[0][2] = 2676ns;
slave_timing[2][96+0].t_rxd2[2][0] = 1656ns;
slave_timing[2][96+0].t_rxd2[1][2] = 2235ns;
slave_timing[2][96+0].t_rxd2[2][1] = 2155ns;

slave_timing[2][96+1].info_corner          = 4;
slave_timing[2][96+1].info_temp__j__       = 125;
slave_timing[2][96+1].info_i__quite_rec__  = 0.006000000;
slave_timing[2][96+1].info_dtr__ib__       = -1;
slave_timing[2][96+1].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+1].info_i__max_slave__  = 0.025000000;
slave_timing[2][96+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][96+1].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+1].t_rxd1[0][1] = 2112ns;
slave_timing[2][96+1].t_rxd1[1][0] = 2232ns;
slave_timing[2][96+1].t_rxd1[0][2] = 1610ns;
slave_timing[2][96+1].t_rxd1[2][0] = 2685ns;
slave_timing[2][96+1].t_rxd2[0][2] = 2517ns;
slave_timing[2][96+1].t_rxd2[2][0] = 1773ns;
slave_timing[2][96+1].t_rxd2[1][2] = 2008ns;
slave_timing[2][96+1].t_rxd2[2][1] = 2394ns;

slave_timing[2][96+2].info_corner          = 4;
slave_timing[2][96+2].info_temp__j__       = 125;
slave_timing[2][96+2].info_i__quite_rec__  = 0.006000000;
slave_timing[2][96+2].info_dtr__ib__       = 1;
slave_timing[2][96+2].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+2].info_i__max_slave__  = 0.023000000;
slave_timing[2][96+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][96+2].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+2].t_rxd1[0][1] = 2217ns;
slave_timing[2][96+2].t_rxd1[1][0] = 2109ns;
slave_timing[2][96+2].t_rxd1[0][2] = 1663ns;
slave_timing[2][96+2].t_rxd1[2][0] = 2586ns;
slave_timing[2][96+2].t_rxd2[0][2] = 2769ns;
slave_timing[2][96+2].t_rxd2[2][0] = 1557ns;
slave_timing[2][96+2].t_rxd2[1][2] = 2397ns;
slave_timing[2][96+2].t_rxd2[2][1] = 1999ns;

slave_timing[2][96+3].info_corner          = 4;
slave_timing[2][96+3].info_temp__j__       = 125;
slave_timing[2][96+3].info_i__quite_rec__  = 0.006000000;
slave_timing[2][96+3].info_dtr__ib__       = 1;
slave_timing[2][96+3].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+3].info_i__max_slave__  = 0.025000000;
slave_timing[2][96+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][96+3].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+3].t_rxd1[0][1] = 2129ns;
slave_timing[2][96+3].t_rxd1[1][0] = 2178ns;
slave_timing[2][96+3].t_rxd1[0][2] = 1614ns;
slave_timing[2][96+3].t_rxd1[2][0] = 2630ns;
slave_timing[2][96+3].t_rxd2[0][2] = 2588ns;
slave_timing[2][96+3].t_rxd2[2][0] = 1691ns;
slave_timing[2][96+3].t_rxd2[1][2] = 2135ns;
slave_timing[2][96+3].t_rxd2[2][1] = 2223ns;

slave_timing[2][96+4].info_corner          = 4;
slave_timing[2][96+4].info_temp__j__       = 125;
slave_timing[2][96+4].info_i__quite_rec__  = 0.006000000;
slave_timing[2][96+4].info_dtr__ib__       = -1;
slave_timing[2][96+4].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+4].info_i__max_slave__  = 0.023000000;
slave_timing[2][96+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][96+4].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+4].t_rxd1[0][1] = 2377ns;
slave_timing[2][96+4].t_rxd1[1][0] = 2307ns;
slave_timing[2][96+4].t_rxd1[0][2] = 1808ns;
slave_timing[2][96+4].t_rxd1[2][0] = 2766ns;
slave_timing[2][96+4].t_rxd2[0][2] = 2703ns;
slave_timing[2][96+4].t_rxd2[2][0] = 1684ns;
slave_timing[2][96+4].t_rxd2[1][2] = 2260ns;
slave_timing[2][96+4].t_rxd2[2][1] = 2184ns;

slave_timing[2][96+5].info_corner          = 4;
slave_timing[2][96+5].info_temp__j__       = 125;
slave_timing[2][96+5].info_i__quite_rec__  = 0.006000000;
slave_timing[2][96+5].info_dtr__ib__       = -1;
slave_timing[2][96+5].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+5].info_i__max_slave__  = 0.025000000;
slave_timing[2][96+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][96+5].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+5].t_rxd1[0][1] = 2284ns;
slave_timing[2][96+5].t_rxd1[1][0] = 2378ns;
slave_timing[2][96+5].t_rxd1[0][2] = 1756ns;
slave_timing[2][96+5].t_rxd1[2][0] = 2809ns;
slave_timing[2][96+5].t_rxd2[0][2] = 2554ns;
slave_timing[2][96+5].t_rxd2[2][0] = 1797ns;
slave_timing[2][96+5].t_rxd2[1][2] = 2033ns;
slave_timing[2][96+5].t_rxd2[2][1] = 2412ns;

slave_timing[2][96+6].info_corner          = 4;
slave_timing[2][96+6].info_temp__j__       = 125;
slave_timing[2][96+6].info_i__quite_rec__  = 0.006000000;
slave_timing[2][96+6].info_dtr__ib__       = 1;
slave_timing[2][96+6].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+6].info_i__max_slave__  = 0.023000000;
slave_timing[2][96+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][96+6].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+6].t_rxd1[0][1] = 2386ns;
slave_timing[2][96+6].t_rxd1[1][0] = 2245ns;
slave_timing[2][96+6].t_rxd1[0][2] = 1808ns;
slave_timing[2][96+6].t_rxd1[2][0] = 2707ns;
slave_timing[2][96+6].t_rxd2[0][2] = 2791ns;
slave_timing[2][96+6].t_rxd2[2][0] = 1583ns;
slave_timing[2][96+6].t_rxd2[1][2] = 2411ns;
slave_timing[2][96+6].t_rxd2[2][1] = 2020ns;

slave_timing[2][96+7].info_corner          = 4;
slave_timing[2][96+7].info_temp__j__       = 125;
slave_timing[2][96+7].info_i__quite_rec__  = 0.006000000;
slave_timing[2][96+7].info_dtr__ib__       = 1;
slave_timing[2][96+7].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+7].info_i__max_slave__  = 0.025000000;
slave_timing[2][96+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][96+7].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+7].t_rxd1[0][1] = 2301ns;
slave_timing[2][96+7].t_rxd1[1][0] = 2294ns;
slave_timing[2][96+7].t_rxd1[0][2] = 1758ns;
slave_timing[2][96+7].t_rxd1[2][0] = 2749ns;
slave_timing[2][96+7].t_rxd2[0][2] = 2618ns;
slave_timing[2][96+7].t_rxd2[2][0] = 1712ns;
slave_timing[2][96+7].t_rxd2[1][2] = 2186ns;
slave_timing[2][96+7].t_rxd2[2][1] = 2215ns;

slave_timing[2][96+8].info_corner          = 4;
slave_timing[2][96+8].info_temp__j__       = 125;
slave_timing[2][96+8].info_i__quite_rec__  = 0.003000000;
slave_timing[2][96+8].info_dtr__ib__       = -1;
slave_timing[2][96+8].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+8].info_i__max_slave__  = 0.023000000;
slave_timing[2][96+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][96+8].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+8].t_rxd1[0][1] = 2166ns;
slave_timing[2][96+8].t_rxd1[1][0] = 2129ns;
slave_timing[2][96+8].t_rxd1[0][2] = 1629ns;
slave_timing[2][96+8].t_rxd1[2][0] = 2588ns;
slave_timing[2][96+8].t_rxd2[0][2] = 2637ns;
slave_timing[2][96+8].t_rxd2[2][0] = 1625ns;
slave_timing[2][96+8].t_rxd2[1][2] = 2215ns;
slave_timing[2][96+8].t_rxd2[2][1] = 2117ns;

slave_timing[2][96+9].info_corner          = 4;
slave_timing[2][96+9].info_temp__j__       = 125;
slave_timing[2][96+9].info_i__quite_rec__  = 0.003000000;
slave_timing[2][96+9].info_dtr__ib__       = -1;
slave_timing[2][96+9].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+9].info_i__max_slave__  = 0.025000000;
slave_timing[2][96+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][96+9].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+9].t_rxd1[0][1] = 2075ns;
slave_timing[2][96+9].t_rxd1[1][0] = 2195ns;
slave_timing[2][96+9].t_rxd1[0][2] = 1581ns;
slave_timing[2][96+9].t_rxd1[2][0] = 2636ns;
slave_timing[2][96+9].t_rxd2[0][2] = 2481ns;
slave_timing[2][96+9].t_rxd2[2][0] = 1742ns;
slave_timing[2][96+9].t_rxd2[1][2] = 1994ns;
slave_timing[2][96+9].t_rxd2[2][1] = 2350ns;

slave_timing[2][96+10].info_corner          = 4;
slave_timing[2][96+10].info_temp__j__       = 125;
slave_timing[2][96+10].info_i__quite_rec__  = 0.003000000;
slave_timing[2][96+10].info_dtr__ib__       = 1;
slave_timing[2][96+10].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+10].info_i__max_slave__  = 0.023000000;
slave_timing[2][96+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][96+10].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+10].t_rxd1[0][1] = 2200ns;
slave_timing[2][96+10].t_rxd1[1][0] = 2080ns;
slave_timing[2][96+10].t_rxd1[0][2] = 1613ns;
slave_timing[2][96+10].t_rxd1[2][0] = 2545ns;
slave_timing[2][96+10].t_rxd2[0][2] = 2707ns;
slave_timing[2][96+10].t_rxd2[2][0] = 1515ns;
slave_timing[2][96+10].t_rxd2[1][2] = 2374ns;
slave_timing[2][96+10].t_rxd2[2][1] = 1939ns;

slave_timing[2][96+11].info_corner          = 4;
slave_timing[2][96+11].info_temp__j__       = 125;
slave_timing[2][96+11].info_i__quite_rec__  = 0.003000000;
slave_timing[2][96+11].info_dtr__ib__       = 1;
slave_timing[2][96+11].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+11].info_i__max_slave__  = 0.025000000;
slave_timing[2][96+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][96+11].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+11].t_rxd1[0][1] = 2122ns;
slave_timing[2][96+11].t_rxd1[1][0] = 2138ns;
slave_timing[2][96+11].t_rxd1[0][2] = 1594ns;
slave_timing[2][96+11].t_rxd1[2][0] = 2589ns;
slave_timing[2][96+11].t_rxd2[0][2] = 2561ns;
slave_timing[2][96+11].t_rxd2[2][0] = 1645ns;
slave_timing[2][96+11].t_rxd2[1][2] = 2113ns;
slave_timing[2][96+11].t_rxd2[2][1] = 2169ns;

slave_timing[2][96+12].info_corner          = 4;
slave_timing[2][96+12].info_temp__j__       = 125;
slave_timing[2][96+12].info_i__quite_rec__  = 0.003000000;
slave_timing[2][96+12].info_dtr__ib__       = -1;
slave_timing[2][96+12].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+12].info_i__max_slave__  = 0.023000000;
slave_timing[2][96+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][96+12].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+12].t_rxd1[0][1] = 2353ns;
slave_timing[2][96+12].t_rxd1[1][0] = 2267ns;
slave_timing[2][96+12].t_rxd1[0][2] = 1793ns;
slave_timing[2][96+12].t_rxd1[2][0] = 2718ns;
slave_timing[2][96+12].t_rxd2[0][2] = 2663ns;
slave_timing[2][96+12].t_rxd2[2][0] = 1649ns;
slave_timing[2][96+12].t_rxd2[1][2] = 2272ns;
slave_timing[2][96+12].t_rxd2[2][1] = 2112ns;

slave_timing[2][96+13].info_corner          = 4;
slave_timing[2][96+13].info_temp__j__       = 125;
slave_timing[2][96+13].info_i__quite_rec__  = 0.003000000;
slave_timing[2][96+13].info_dtr__ib__       = -1;
slave_timing[2][96+13].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+13].info_i__max_slave__  = 0.025000000;
slave_timing[2][96+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][96+13].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+13].t_rxd1[0][1] = 2269ns;
slave_timing[2][96+13].t_rxd1[1][0] = 2348ns;
slave_timing[2][96+13].t_rxd1[0][2] = 1742ns;
slave_timing[2][96+13].t_rxd1[2][0] = 2762ns;
slave_timing[2][96+13].t_rxd2[0][2] = 2515ns;
slave_timing[2][96+13].t_rxd2[2][0] = 1767ns;
slave_timing[2][96+13].t_rxd2[1][2] = 2008ns;
slave_timing[2][96+13].t_rxd2[2][1] = 2364ns;

slave_timing[2][96+14].info_corner          = 4;
slave_timing[2][96+14].info_temp__j__       = 125;
slave_timing[2][96+14].info_i__quite_rec__  = 0.003000000;
slave_timing[2][96+14].info_dtr__ib__       = 1;
slave_timing[2][96+14].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+14].info_i__max_slave__  = 0.023000000;
slave_timing[2][96+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][96+14].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+14].t_rxd1[0][1] = 2386ns;
slave_timing[2][96+14].t_rxd1[1][0] = 2223ns;
slave_timing[2][96+14].t_rxd1[0][2] = 1798ns;
slave_timing[2][96+14].t_rxd1[2][0] = 2660ns;
slave_timing[2][96+14].t_rxd2[0][2] = 2753ns;
slave_timing[2][96+14].t_rxd2[2][0] = 1539ns;
slave_timing[2][96+14].t_rxd2[1][2] = 2387ns;
slave_timing[2][96+14].t_rxd2[2][1] = 1967ns;

slave_timing[2][96+15].info_corner          = 4;
slave_timing[2][96+15].info_temp__j__       = 125;
slave_timing[2][96+15].info_i__quite_rec__  = 0.003000000;
slave_timing[2][96+15].info_dtr__ib__       = 1;
slave_timing[2][96+15].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+15].info_i__max_slave__  = 0.025000000;
slave_timing[2][96+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][96+15].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+15].t_rxd1[0][1] = 2298ns;
slave_timing[2][96+15].t_rxd1[1][0] = 2261ns;
slave_timing[2][96+15].t_rxd1[0][2] = 1750ns;
slave_timing[2][96+15].t_rxd1[2][0] = 2709ns;
slave_timing[2][96+15].t_rxd2[0][2] = 2581ns;
slave_timing[2][96+15].t_rxd2[2][0] = 1669ns;
slave_timing[2][96+15].t_rxd2[1][2] = 2137ns;
slave_timing[2][96+15].t_rxd2[2][1] = 2190ns;

slave_timing[2][96+16].info_corner          = 4;
slave_timing[2][96+16].info_temp__j__       = 125;
slave_timing[2][96+16].info_i__quite_rec__  = 0.000000000;
slave_timing[2][96+16].info_dtr__ib__       = -1;
slave_timing[2][96+16].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+16].info_i__max_slave__  = 0.023000000;
slave_timing[2][96+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][96+16].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+16].t_rxd1[0][1] = 2148ns;
slave_timing[2][96+16].t_rxd1[1][0] = 2104ns;
slave_timing[2][96+16].t_rxd1[0][2] = 1611ns;
slave_timing[2][96+16].t_rxd1[2][0] = 2552ns;
slave_timing[2][96+16].t_rxd2[0][2] = 2596ns;
slave_timing[2][96+16].t_rxd2[2][0] = 1585ns;
slave_timing[2][96+16].t_rxd2[1][2] = 2191ns;
slave_timing[2][96+16].t_rxd2[2][1] = 2071ns;

slave_timing[2][96+17].info_corner          = 4;
slave_timing[2][96+17].info_temp__j__       = 125;
slave_timing[2][96+17].info_i__quite_rec__  = 0.000000000;
slave_timing[2][96+17].info_dtr__ib__       = -1;
slave_timing[2][96+17].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+17].info_i__max_slave__  = 0.025000000;
slave_timing[2][96+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][96+17].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+17].t_rxd1[0][1] = 2048ns;
slave_timing[2][96+17].t_rxd1[1][0] = 2164ns;
slave_timing[2][96+17].t_rxd1[0][2] = 1565ns;
slave_timing[2][96+17].t_rxd1[2][0] = 2593ns;
slave_timing[2][96+17].t_rxd2[0][2] = 2442ns;
slave_timing[2][96+17].t_rxd2[2][0] = 1703ns;
slave_timing[2][96+17].t_rxd2[1][2] = 1963ns;
slave_timing[2][96+17].t_rxd2[2][1] = 2287ns;

slave_timing[2][96+18].info_corner          = 4;
slave_timing[2][96+18].info_temp__j__       = 125;
slave_timing[2][96+18].info_i__quite_rec__  = 0.000000000;
slave_timing[2][96+18].info_dtr__ib__       = 1;
slave_timing[2][96+18].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+18].info_i__max_slave__  = 0.023000000;
slave_timing[2][96+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][96+18].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+18].t_rxd1[0][1] = 2172ns;
slave_timing[2][96+18].t_rxd1[1][0] = 2050ns;
slave_timing[2][96+18].t_rxd1[0][2] = 1620ns;
slave_timing[2][96+18].t_rxd1[2][0] = 2512ns;
slave_timing[2][96+18].t_rxd2[0][2] = 2694ns;
slave_timing[2][96+18].t_rxd2[2][0] = 1462ns;
slave_timing[2][96+18].t_rxd2[1][2] = 2333ns;
slave_timing[2][96+18].t_rxd2[2][1] = 1896ns;

slave_timing[2][96+19].info_corner          = 4;
slave_timing[2][96+19].info_temp__j__       = 125;
slave_timing[2][96+19].info_i__quite_rec__  = 0.000000000;
slave_timing[2][96+19].info_dtr__ib__       = 1;
slave_timing[2][96+19].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+19].info_i__max_slave__  = 0.025000000;
slave_timing[2][96+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][96+19].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+19].t_rxd1[0][1] = 2074ns;
slave_timing[2][96+19].t_rxd1[1][0] = 2125ns;
slave_timing[2][96+19].t_rxd1[0][2] = 1569ns;
slave_timing[2][96+19].t_rxd1[2][0] = 2552ns;
slave_timing[2][96+19].t_rxd2[0][2] = 2515ns;
slave_timing[2][96+19].t_rxd2[2][0] = 1614ns;
slave_timing[2][96+19].t_rxd2[1][2] = 2084ns;
slave_timing[2][96+19].t_rxd2[2][1] = 2130ns;

slave_timing[2][96+20].info_corner          = 4;
slave_timing[2][96+20].info_temp__j__       = 125;
slave_timing[2][96+20].info_i__quite_rec__  = 0.000000000;
slave_timing[2][96+20].info_dtr__ib__       = -1;
slave_timing[2][96+20].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+20].info_i__max_slave__  = 0.023000000;
slave_timing[2][96+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][96+20].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+20].t_rxd1[0][1] = 2357ns;
slave_timing[2][96+20].t_rxd1[1][0] = 2246ns;
slave_timing[2][96+20].t_rxd1[0][2] = 1793ns;
slave_timing[2][96+20].t_rxd1[2][0] = 2670ns;
slave_timing[2][96+20].t_rxd2[0][2] = 2611ns;
slave_timing[2][96+20].t_rxd2[2][0] = 1601ns;
slave_timing[2][96+20].t_rxd2[1][2] = 2245ns;
slave_timing[2][96+20].t_rxd2[2][1] = 2058ns;

slave_timing[2][96+21].info_corner          = 4;
slave_timing[2][96+21].info_temp__j__       = 125;
slave_timing[2][96+21].info_i__quite_rec__  = 0.000000000;
slave_timing[2][96+21].info_dtr__ib__       = -1;
slave_timing[2][96+21].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+21].info_i__max_slave__  = 0.025000000;
slave_timing[2][96+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][96+21].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+21].t_rxd1[0][1] = 2265ns;
slave_timing[2][96+21].t_rxd1[1][0] = 2307ns;
slave_timing[2][96+21].t_rxd1[0][2] = 1743ns;
slave_timing[2][96+21].t_rxd1[2][0] = 2720ns;
slave_timing[2][96+21].t_rxd2[0][2] = 2465ns;
slave_timing[2][96+21].t_rxd2[2][0] = 1727ns;
slave_timing[2][96+21].t_rxd2[1][2] = 2015ns;
slave_timing[2][96+21].t_rxd2[2][1] = 2280ns;

slave_timing[2][96+22].info_corner          = 4;
slave_timing[2][96+22].info_temp__j__       = 125;
slave_timing[2][96+22].info_i__quite_rec__  = 0.000000000;
slave_timing[2][96+22].info_dtr__ib__       = 1;
slave_timing[2][96+22].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+22].info_i__max_slave__  = 0.023000000;
slave_timing[2][96+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][96+22].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+22].t_rxd1[0][1] = 2371ns;
slave_timing[2][96+22].t_rxd1[1][0] = 2188ns;
slave_timing[2][96+22].t_rxd1[0][2] = 1797ns;
slave_timing[2][96+22].t_rxd1[2][0] = 2629ns;
slave_timing[2][96+22].t_rxd2[0][2] = 2703ns;
slave_timing[2][96+22].t_rxd2[2][0] = 1478ns;
slave_timing[2][96+22].t_rxd2[1][2] = 2345ns;
slave_timing[2][96+22].t_rxd2[2][1] = 1901ns;

slave_timing[2][96+23].info_corner          = 4;
slave_timing[2][96+23].info_temp__j__       = 125;
slave_timing[2][96+23].info_i__quite_rec__  = 0.000000000;
slave_timing[2][96+23].info_dtr__ib__       = 1;
slave_timing[2][96+23].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+23].info_i__max_slave__  = 0.025000000;
slave_timing[2][96+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][96+23].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+23].t_rxd1[0][1] = 2288ns;
slave_timing[2][96+23].t_rxd1[1][0] = 2254ns;
slave_timing[2][96+23].t_rxd1[0][2] = 1747ns;
slave_timing[2][96+23].t_rxd1[2][0] = 2673ns;
slave_timing[2][96+23].t_rxd2[0][2] = 2536ns;
slave_timing[2][96+23].t_rxd2[2][0] = 1632ns;
slave_timing[2][96+23].t_rxd2[1][2] = 2113ns;
slave_timing[2][96+23].t_rxd2[2][1] = 2142ns;

slave_timing[2][96+24].info_corner          = 4;
slave_timing[2][96+24].info_temp__j__       = 125;
slave_timing[2][96+24].info_i__quite_rec__  = 0.040000000;
slave_timing[2][96+24].info_dtr__ib__       = -1;
slave_timing[2][96+24].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+24].info_i__max_slave__  = 0.023000000;
slave_timing[2][96+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][96+24].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+24].t_rxd1[0][1] = 2251ns;
slave_timing[2][96+24].t_rxd1[1][0] = 2225ns;
slave_timing[2][96+24].t_rxd1[0][2] = 1729ns;
slave_timing[2][96+24].t_rxd1[2][0] = 2754ns;
slave_timing[2][96+24].t_rxd2[0][2] = 2958ns;
slave_timing[2][96+24].t_rxd2[2][0] = 1870ns;
slave_timing[2][96+24].t_rxd2[1][2] = 2494ns;
slave_timing[2][96+24].t_rxd2[2][1] = 2438ns;

slave_timing[2][96+25].info_corner          = 4;
slave_timing[2][96+25].info_temp__j__       = 125;
slave_timing[2][96+25].info_i__quite_rec__  = 0.040000000;
slave_timing[2][96+25].info_dtr__ib__       = -1;
slave_timing[2][96+25].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+25].info_i__max_slave__  = 0.025000000;
slave_timing[2][96+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][96+25].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+25].t_rxd1[0][1] = 2173ns;
slave_timing[2][96+25].t_rxd1[1][0] = 2306ns;
slave_timing[2][96+25].t_rxd1[0][2] = 1681ns;
slave_timing[2][96+25].t_rxd1[2][0] = 2803ns;
slave_timing[2][96+25].t_rxd2[0][2] = 2792ns;
slave_timing[2][96+25].t_rxd2[2][0] = 1993ns;
slave_timing[2][96+25].t_rxd2[1][2] = 2271ns;
slave_timing[2][96+25].t_rxd2[2][1] = 2639ns;

slave_timing[2][96+26].info_corner          = 4;
slave_timing[2][96+26].info_temp__j__       = 125;
slave_timing[2][96+26].info_i__quite_rec__  = 0.040000000;
slave_timing[2][96+26].info_dtr__ib__       = 1;
slave_timing[2][96+26].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+26].info_i__max_slave__  = 0.023000000;
slave_timing[2][96+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][96+26].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+26].t_rxd1[0][1] = 2319ns;
slave_timing[2][96+26].t_rxd1[1][0] = 2169ns;
slave_timing[2][96+26].t_rxd1[0][2] = 1756ns;
slave_timing[2][96+26].t_rxd1[2][0] = 2711ns;
slave_timing[2][96+26].t_rxd2[0][2] = 3094ns;
slave_timing[2][96+26].t_rxd2[2][0] = 1767ns;
slave_timing[2][96+26].t_rxd2[1][2] = 2688ns;
slave_timing[2][96+26].t_rxd2[2][1] = 2255ns;

slave_timing[2][96+27].info_corner          = 4;
slave_timing[2][96+27].info_temp__j__       = 125;
slave_timing[2][96+27].info_i__quite_rec__  = 0.040000000;
slave_timing[2][96+27].info_dtr__ib__       = 1;
slave_timing[2][96+27].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+27].info_i__max_slave__  = 0.025000000;
slave_timing[2][96+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][96+27].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+27].t_rxd1[0][1] = 2236ns;
slave_timing[2][96+27].t_rxd1[1][0] = 2249ns;
slave_timing[2][96+27].t_rxd1[0][2] = 1718ns;
slave_timing[2][96+27].t_rxd1[2][0] = 2769ns;
slave_timing[2][96+27].t_rxd2[0][2] = 2900ns;
slave_timing[2][96+27].t_rxd2[2][0] = 1905ns;
slave_timing[2][96+27].t_rxd2[1][2] = 2410ns;
slave_timing[2][96+27].t_rxd2[2][1] = 2491ns;

slave_timing[2][96+28].info_corner          = 4;
slave_timing[2][96+28].info_temp__j__       = 125;
slave_timing[2][96+28].info_i__quite_rec__  = 0.040000000;
slave_timing[2][96+28].info_dtr__ib__       = -1;
slave_timing[2][96+28].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+28].info_i__max_slave__  = 0.023000000;
slave_timing[2][96+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][96+28].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+28].t_rxd1[0][1] = 2332ns;
slave_timing[2][96+28].t_rxd1[1][0] = 2638ns;
slave_timing[2][96+28].t_rxd1[0][2] = 1815ns;
slave_timing[2][96+28].t_rxd1[2][0] = 3568ns;
slave_timing[2][96+28].t_rxd2[0][2] = 3879ns;
slave_timing[2][96+28].t_rxd2[2][0] = 2446ns;
slave_timing[2][96+28].t_rxd2[1][2] = 3324ns;
slave_timing[2][96+28].t_rxd2[2][1] = 3263ns;

slave_timing[2][96+29].info_corner          = 4;
slave_timing[2][96+29].info_temp__j__       = 125;
slave_timing[2][96+29].info_i__quite_rec__  = 0.040000000;
slave_timing[2][96+29].info_dtr__ib__       = -1;
slave_timing[2][96+29].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+29].info_i__max_slave__  = 0.025000000;
slave_timing[2][96+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][96+29].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+29].t_rxd1[0][1] = 2256ns;
slave_timing[2][96+29].t_rxd1[1][0] = 2749ns;
slave_timing[2][96+29].t_rxd1[0][2] = 1785ns;
slave_timing[2][96+29].t_rxd1[2][0] = 3678ns;
slave_timing[2][96+29].t_rxd2[0][2] = 3596ns;
slave_timing[2][96+29].t_rxd2[2][0] = 2617ns;
slave_timing[2][96+29].t_rxd2[1][2] = 2943ns;
slave_timing[2][96+29].t_rxd2[2][1] = 3673ns;

slave_timing[2][96+30].info_corner          = 4;
slave_timing[2][96+30].info_temp__j__       = 125;
slave_timing[2][96+30].info_i__quite_rec__  = 0.040000000;
slave_timing[2][96+30].info_dtr__ib__       = 1;
slave_timing[2][96+30].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+30].info_i__max_slave__  = 0.023000000;
slave_timing[2][96+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][96+30].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+30].t_rxd1[0][1] = 2395ns;
slave_timing[2][96+30].t_rxd1[1][0] = 2494ns;
slave_timing[2][96+30].t_rxd1[0][2] = 1862ns;
slave_timing[2][96+30].t_rxd1[2][0] = 3446ns;
slave_timing[2][96+30].t_rxd2[0][2] = 4131ns;
slave_timing[2][96+30].t_rxd2[2][0] = 2300ns;
slave_timing[2][96+30].t_rxd2[1][2] = 3629ns;
slave_timing[2][96+30].t_rxd2[2][1] = 2987ns;

slave_timing[2][96+31].info_corner          = 4;
slave_timing[2][96+31].info_temp__j__       = 125;
slave_timing[2][96+31].info_i__quite_rec__  = 0.040000000;
slave_timing[2][96+31].info_dtr__ib__       = 1;
slave_timing[2][96+31].info_i__offset_rec__ = 0.000000000;
slave_timing[2][96+31].info_i__max_slave__  = 0.025000000;
slave_timing[2][96+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][96+31].info_r__dsi_bus__    = 5.000;

slave_timing[2][96+31].t_rxd1[0][1] = 2305ns;
slave_timing[2][96+31].t_rxd1[1][0] = 2630ns;
slave_timing[2][96+31].t_rxd1[0][2] = 1816ns;
slave_timing[2][96+31].t_rxd1[2][0] = 3553ns;
slave_timing[2][96+31].t_rxd2[0][2] = 3768ns;
slave_timing[2][96+31].t_rxd2[2][0] = 2488ns;
slave_timing[2][96+31].t_rxd2[1][2] = 3186ns;
slave_timing[2][96+31].t_rxd2[2][1] = 3357ns;

/**
 * Package: unit_test_pkg
 * 
 * package for unit testing
 */
package unit_test_pkg;
	import uvm_pkg::*;
	import common_pkg::*;
	import common_env_pkg::*;
	import spi_pkg::*;
	import dsi3_slave_pkg::*;
	import dsi3_pkg::*;
	import project_pkg::*;
	import common_test_pkg::*;
	import digital_signal_pkg::*;
	import regmodel_pkg::*;
	
	`include "dsi3_master_configuration_listener.svh"
	
	`uvm_analysis_imp_decl(_buffer_writer)
	`uvm_analysis_imp_decl(_elip_writer)
	`uvm_analysis_imp_decl(_frame_writer)
	
	`include "default_comparer.svh"
	
	`include "dsi3_slave_test_driver.svh"
	`include "dsi3_receiver_test_slave_sequence.svh"
	`include "receive_service.svh"
	
	`include "m52142b_slave_timing.svh"
	
	`include "top_config.svh"
	`include "top_env.svh"
	`include "top_test.svh"
	`include "chip_time_iterator.svh"

endpackage




`include "sub_sequences/pdcm/upload_tdma_scheme_seq.svh"
`include "sub_sequences/pdcm/upload_random_valid_tdma_schemes_seq.svh"
`include "sub_sequences/pdcm/upload_random_invalid_tdma_schemes_seq.svh"
`include "sub_sequences/pdcm/upload_tdma_scheme_and_start_pdcm_in_one_frame_seq.svh"
`include "sub_sequences/pdcm/start_pdcm_without_valid_tdma_scheme_seq.svh"
`include "sub_sequences/pdcm/single_pdcm_on_all_channels_seq.svh"
`include "sub_sequences/pdcm/single_pdcm_on_all_channels_fail_seq.svh"
`include "sub_sequences/pdcm/single_pdcm_on_single_channel_seq.svh"
`include "sub_sequences/pdcm/pdcm_early_single_packet_seq.svh"
`include "sub_sequences/pdcm/pdcm_late_single_packet_seq.svh"
`include "sub_sequences/pdcm/pdcm_packet_count_error_seq.svh"
`include "sub_sequences/pdcm/pdcm_maximum_packet_count_error_seq.svh"
`include "sub_sequences/pdcm/pdcm_symbol_count_error_seq.svh"
`include "sub_sequences/pdcm/pdcm_symbol_coding_error_seq.svh"
`include "sub_sequences/pdcm/pdcm_voltage_error_seq.svh"
`include "sub_sequences/pdcm/pdcm_voltage_error_before_slave_answer_seq.svh"
`include "sub_sequences/pdcm/pdcm_clock_ref_error_seq.svh"
`include "sub_sequences/pdcm/pdcm_clock_ref_error_during_pdcm_pulse_transmission_seq.svh"
`include "sub_sequences/pdcm/pdcm_receive_packet_with_more_than_255_symbols_seq.svh"
`include "sub_sequences/pdcm/pdcm_with_maximum_pulse_count_seq.svh"
`include "sub_sequences/pdcm/pdcm_min_max_periods_seq.svh"
`include "sub_sequences/pdcm/pdcm_packet_start_before_t__PDCM_START__seq.svh"
`include "sub_sequences/pdcm/pdcm_packets_too_late_seq.svh"
`include "sub_sequences/pdcm/pdcm_symbol_noise_on_all_channels_seq.svh"
`include "sub_sequences/pdcm/pdcm_chip_noise_on_all_channels_seq.svh"
`include "sub_sequences/pdcm/pdcm_single_packet_split_by_end_of_period_seq.svh"
`include "sub_sequences/pdcm/pdcm_short_inter_packet_gaps_seq.svh"
`include "sub_sequences/pdcm/pdcm_long_packets_end_at_receive_timeout_seq.svh"
`include "sub_sequences/pdcm/pdcm_ram_burst_read_seq.svh"
`include "sub_sequences/pdcm/pdcm_fill_buffer_seq.svh"
`include "sub_sequences/pdcm/pdcm_denso_one_missing_and_one_too_large_packet_seq.svh"
`include "sub_sequences/pdcm/pdcm_denso_one_moving_packet_seq.svh"
`include "sub_sequences/pdcm/pdcm_random_denso_scheme_on_all_channels_seq.svh"
`include "sub_sequences/pdcm/pdcm_random_denso_15_scheme_on_all_channels_seq.svh"
`include "sub_sequences/pdcm/pdcm_denso_scheme_all_source_ids_seq.svh"
`include "sub_sequences/pdcm/pdcm_measure_t__PDCM_END__seq.svh"

`include "sub_sequences/pdcm/pdcm_denso_15_single_missing_packet_seq.svh"
`include "sub_sequences/pdcm/pdcm_denso_15_random_missing_packets_seq.svh"
`include "sub_sequences/pdcm/pdcm_read_all_packets_missing_seq.svh"
`include "sub_sequences/pdcm/pdcm_read_empty_data_seq.svh"
`include "sub_sequences/pdcm/pdcm_read_without_pdcm_on_one_channel_scheme_seq.svh"
`include "sub_sequences/pdcm/pdcm_read_without_pdcm_scheme_seq.svh"

`include "sub_sequences/pdcm/random_pdcm_and_different_bit_chip_times_seq.svh"
`include "sub_sequences/pdcm/random_pdcm_and_read_data_seq.svh"
`include "sub_sequences/pdcm/random_pdcm_and_read_multiple_packets_seq.svh"
`include "sub_sequences/pdcm/random_pdcm_fill_data_buffer_seq.svh"
`include "sub_sequences/pdcm/random_pdcm_seq.svh"

`include "sub_sequences/crm/crm_single_channel_transmit_seq.svh"
`include "sub_sequences/crm/crm_many_on_one_channel_one_on_all_channels_seq.svh"
`include "sub_sequences/crm/crm_read_data_using_multiple_tx_crc_seq.svh"
`include "sub_sequences/crm/crm_without_slave_answer_seq.svh"
`include "sub_sequences/crm/crm_transmit_and_read_in_one_frame_seq.svh"
`include "sub_sequences/crm/crm_many_crm_in_one_spi_frame_started_with_tx_crc_seq.svh"
`include "sub_sequences/crm/crm_wrong_symbol_counts_seq.svh"
`include "sub_sequences/crm/crm_late_long_slave_answers_seq.svh"
`include "sub_sequences/crm/crm_late_short_slave_answers_seq.svh"
`include "sub_sequences/crm/crm_very_long_slave_answers_seq.svh"
`include "sub_sequences/crm/crm_very_long_slave_answers_with_additional_crm_seq.svh"
`include "sub_sequences/crm/crm_two_short_slave_answers_seq.svh"
`include "sub_sequences/crm/crm_clock_ref_error_during_crm_transmission_seq.svh"
`include "sub_sequences/crm/crm_clock_ref_error_in_crm_for_all_channels_seq.svh"
`include "sub_sequences/crm/crm_clock_ref_inside_crm_transmission_seq.svh"
`include "sub_sequences/crm/crm_clock_ref_disable_during_crm_transmission_seq.svh"
`include "sub_sequences/crm/crm_clock_ref_error_during_crm_transmission_without_slave_answer_seq.svh"
`include "sub_sequences/crm/crm_voltage_error_in_crm_for_all_channels_seq.svh"
`include "sub_sequences/crm/crm_symbol_coding_error_in_crm_for_all_channels_seq.svh"
`include "sub_sequences/crm/crm_chip_coding_error_in_crm_for_all_channels_seq.svh"
`include "sub_sequences/crm/crm_crc_en_seq.svh"
`include "sub_sequences/crm/crm_multiple_crms_in_one_command_frame_seq.svh"
`include "sub_sequences/crm/crm_multiple_broadcast_crms_in_one_command_frame_seq.svh"
`include "sub_sequences/crm/crm_symbol_noise_on_all_channels_seq.svh"
`include "sub_sequences/crm/crm_dsi_fast_config_access_seq.svh"
`include "sub_sequences/crm/crm_check_different_chiptimes_and_bittimes_seq.svh"
`include "sub_sequences/crm/crm_fill_buffer_seq.svh"
`include "sub_sequences/crm/crm_random_on_different_channels_seq.svh"
`include "sub_sequences/crm/crm_disable_clock_ref_during_transmission_p52143_697_seq.svh"
`include "sub_sequences/crm/crm_read_empty_data_seq.svh"
`include "sub_sequences/crm/crm_CRM_TIME_lower_than_transmission_time_seq.svh"
`include "sub_sequences/crm/crm_CRM_TIME_NR_lower_than_transmission_time_seq.svh"
`include "sub_sequences/crm/crm_maximum_CRM_TIME_seq.svh"
`include "sub_sequences/crm/crm_maximum_CRM_TIME_NR_seq.svh"
`include "sub_sequences/crm/crm_maximum_CRM_TIME_with_multiple_answers_seq.svh"
`include "sub_sequences/crm/crm_CRM_TIME_change_during_crm_transmission_seq.svh"
`include "sub_sequences/crm/crm_read_status_during_reception_seq.svh"
`include "sub_sequences/crm/crm_with_ffff_data_seq.svh"

`include "sub_sequences/discovery/dsi3_random_discovery_mode_seq.svh"
`include "sub_sequences/discovery/dsi3_discovery_mode_without_slaves_seq.svh"
`include "sub_sequences/discovery/dsi3_discovery_mode_overflow_seq.svh"

`include "sub_sequences/register/register_check_ic_revision_seq.svh"
`include "sub_sequences/register/register_read_tb_cnt_register_seq.svh"
`include "sub_sequences/register/register_check_ring_buffers_seq.svh"
`include "sub_sequences/register/register_miso_crc_example_seq.svh"
`include "sub_sequences/register/register_irq_en_enable_all_irqs_seq.svh"
`include "sub_sequences/register/register_dsi_irq_en_frontdoor_access_seq.svh"
`include "sub_sequences/register/register_multiple_writes_in_one_frame_seq.svh"
`include "sub_sequences/register/register_multiple_writes_with_tx_crc_in_one_frame_seq.svh"
`include "sub_sequences/register/register_multiple_writes_with_tx_crc_in_one_wrong_crc_frame_seq.svh"
`include "sub_sequences/register/register_write_to_invalid_addresses_seq.svh"
`include "sub_sequences/register/register_spi_burst_read_to_improve_coverage_seq.svh"
`include "sub_sequences/register/register_spi_burst_read_zero_address_seq.svh"
`include "sub_sequences/register/register_jtag_burst_read_to_improve_coverage_seq.svh"
`include "sub_sequences/register/register_read_ic_revision_during_startup_seq.svh"

`include "sub_sequences/spec/spec_Sync_CRM_on_DSI_seq.sv"
`include "sub_sequences/spec/spec_Sync_IDLE_DSI_seq.sv"
`include "sub_sequences/spec/spec_CRM_command_seq.sv"
`include "sub_sequences/spec/spec_CRM_configuration_seq.sv"
`include "sub_sequences/spec/spec_DSI_wait_seq.sv"
`include "sub_sequences/spec/spec_single_frame_pdcm_read_seq.sv"
`include "sub_sequences/spec/spec_multiple_frame_pdcm_read_seq.sv"
`include "sub_sequences/spec/spec_multiple_frame_pdcm_lang_packet_read_seq.sv"
`include "sub_sequences/spec/spec_measurement_command_stack_seq.sv"
`include "sub_sequences/spec/spec_external_Sync_on_DSI_seq.sv"

`include "sub_sequences/spi/spi_access_irq_en_wrong_crc_seq.svh"
`include "sub_sequences/spi/spi_access_irq_en_wrong_and_correct_tx_crc_seq.svh"
`include "sub_sequences/spi/spi_access_irq_en_correct_and_wrong_tx_crc_seq.svh"
`include "sub_sequences/spi/spi_start_frame_with_tx_crc_seq.svh"
`include "sub_sequences/spi/spi_bit_count_errors_seq.svh"
`include "sub_sequences/spi/spi_crc_ends_with_zeros_seq.svh"
`include "sub_sequences/spi/spi_frame_ends_with_reset_command_seq.svh"
`include "sub_sequences/spi/spi_frame_starts_with_reset_command_seq.svh"
`include "sub_sequences/spi/spi_multiple_reset_commands_seq.svh"
`include "sub_sequences/spi/spi_reset_random_command_frame_seq.svh"
`include "sub_sequences/spi/spi_reset_after_valid_command_frame_seq.svh"
`include "sub_sequences/spi/spi_reset_with_bit_count_errors_seq.svh"
`include "sub_sequences/spi/spi_reset_full_spi_command_buffer_seq.svh"
`include "sub_sequences/spi/spi_traffic_with_csb_high_seq.svh"
`include "sub_sequences/spi/spi_incomplete_register_reads_seq.svh"
`include "sub_sequences/spi/spi_incomplete_burst_register_reads_seq.svh"
`include "sub_sequences/spi/spi_incomplete_read_crm_data_seq.svh"
`include "sub_sequences/spi/spi_incomplete_read_crm_data_bit_count_seq.svh"
`include "sub_sequences/spi/spi_incomplete_read_pdcm_denso_15_seq.svh"
`include "sub_sequences/spi/spi_incomplete_read_pdcm_single_packet_seq.svh"
`include "sub_sequences/spi/spi_incomplete_read_pdcm_with_maximum_size_scheme_seq.svh"
`include "sub_sequences/spi/spi_incomplete_reset_command_seq.svh"
`include "sub_sequences/spi/spi_burst_read_with_wrong_tx_crc_seq.svh"
`include "sub_sequences/spi/spi_read_register_and_crm_transmit_with_crc_command_seq.svh"
`include "sub_sequences/spi/spi_hw_fail_during_spi_frame_seq.svh"
`include "sub_sequences/spi/spi_single_command_ignored_seq.svh"
`include "sub_sequences/spi/spi_multiple_command_ignored_seq.svh"

`include "sub_sequences/otp/base_otp_seq.svh"
`include "sub_sequences/otp/otp_random_trimming_seq.svh"
`include "sub_sequences/otp/otp_write_to_ram_seq.svh"
`include "sub_sequences/otp/otp_single_bit_ecc_failure_seq.svh"
`include "sub_sequences/otp/otp_double_bit_ecc_failure_seq.svh"
`include "sub_sequences/otp/otp_mixed_bit_ecc_failure_seq.svh"
`include "sub_sequences/otp/otp_applicative_readout_seq.svh"
`include "sub_sequences/otp/otp_applicative_readout_too_early_seq.svh"
`include "sub_sequences/otp/otp_applicative_readout_much_too_early_seq.svh"
`include "sub_sequences/otp/otp_applicative_readout_fail_by_vcc_vrr_seq.svh"
`include "sub_sequences/otp/otp_applicative_readout_multiple_read_of_same_address_seq.svh"
`include "sub_sequences/otp/otp_applicative_readout_fail_by_vcc_while_reading_seq.svh"
`include "sub_sequences/otp/otp_vcc_uv_during_read_seq.svh"

`include "sub_sequences/debounce/debounce_measure_seq.svh"
`include "sub_sequences/debounce/resb_debounce_measure_seq.svh"
`include "sub_sequences/debounce/vccuv_debounce_measure_seq.svh"
`include "sub_sequences/debounce/ref_fail_debounce_measure_seq.svh"
`include "sub_sequences/debounce/ldo_uv_debounce_measure_seq.svh"
`include "sub_sequences/debounce/ot_debounce_measure_seq.svh"
`include "sub_sequences/debounce/dsi_mon_to_debounce_measure_seq.svh"
`include "sub_sequences/debounce/dsi_uv_debounce_measure_seq.svh"

`include "sub_sequences/jtag/jtag_read_chip_id_seq.svh"

`include "sub_sequences/crm/crm_command_without_data_seq.svh"
`include "sub_sequences/crm/crm_broadcast_and_read_seq.svh"
`include "sub_sequences/crm/single_crm_on_all_channels_seq.svh"
`include "sub_sequences/crm/single_crm_on_all_channels_fail_seq.svh"
`include "sub_sequences/crm/single_crm_on_each_channel_seq.svh"

`include "sub_sequences/wait/base_wait_seq.svh"
`include "sub_sequences/wait/chained_wait_on_each_channel_seq.svh"
`include "sub_sequences/wait/check_wait_register_seq.svh"
`include "sub_sequences/wait/wait_maximum_on_all_channel_seq.svh"
`include "sub_sequences/wait/wait_on_each_channel_seq.svh"

`include "sub_sequences/stop/stop_command_queue_within_command_frame_seq.svh"
`include "sub_sequences/stop/stop_single_pdcm_of_all_channels_seq.svh"
`include "sub_sequences/stop/stop_crm_directly_after_start_seq.svh"
`include "sub_sequences/stop/stop_finite_pdcm_at_random_time_seq.svh"
`include "sub_sequences/stop/stop_infinite_pdcm_at_random_time_seq.svh"
`include "sub_sequences/stop/stop_queued_crm_commands_seq.svh"
`include "sub_sequences/stop/stop_random_command_queue_seq.svh"
`include "sub_sequences/stop/stop_wait_command_seq.svh"

`include "sub_sequences/clear/clear_buffer_and_read_in_one_frame_seq.svh"
`include "sub_sequences/clear/clear_buffer_during_crm_seq.svh"
`include "sub_sequences/clear/clear_buffer_during_pdcm_seq.svh"
`include "sub_sequences/clear/clear_buffer_during_pdcm_fine_delayed_seq.svh"
`include "sub_sequences/clear/clear_crm_and_pdcm_data_buffer_seq.svh"
`include "sub_sequences/clear/clear_crm_data_buffer_seq.svh"
`include "sub_sequences/clear/clear_full_pdcm_buffer_seq.svh"
`include "sub_sequences/clear/clear_pdcm_data_buffer_seq.svh"
`include "sub_sequences/clear/clear_pdcm_data_with_tdma_scheme_upload_seq.svh"
`include "sub_sequences/clear/clear_pdcm_data_with_upload_tdma_packet_seq.svh"
`include "sub_sequences/clear/clear_single_channel_buffer_during_pdcm_seq.svh"

`include "sub_sequences/sync/dsi3_sync_base_seq.sv"
`include "sub_sequences/sync/check_sync_reg_for_crm_seq.svh"
`include "sub_sequences/sync/check_sync_reg_for_pdcm_seq.svh"
`include "sub_sequences/sync/check_sync_reg_for_channel_pairs_seq.svh"
`include "sub_sequences/sync/clear_queue_during_sync_seq.svh"
`include "sub_sequences/sync/clear_queue_of_all_channels_during_sync_seq.svh"
`include "sub_sequences/sync/double_sync_crm_in_different_frames_seq.svh"
`include "sub_sequences/sync/first_sync_at_all_channels_then_single_crms_seq.svh"
`include "sub_sequences/sync/shut_off_during_sync_seq.svh"
`include "sub_sequences/sync/shut_off_before_sync_seq.svh"
`include "sub_sequences/sync/sync_crm_seq.svh"
`include "sub_sequences/sync/sync_multiple_crm_in_different_frames_seq.svh"
`include "sub_sequences/sync/sync_multiple_crm_in_one_frame_seq.svh"
`include "sub_sequences/sync/sync_multiple_crm_per_channel_in_different_frames_seq.svh"
`include "sub_sequences/sync/sync_pdcm_at_all_channels_seq.svh"
`include "sub_sequences/sync/sync_pdcm_seq.svh"
`include "sub_sequences/sync/sync_random_commands_seq.svh"
`include "sub_sequences/sync/wait_for_sync_flag_seq.svh"

`include "sub_sequences/sync_pin/external_sync_crm_seq.svh"
`include "sub_sequences/sync_pin/external_sync_crm_short_pulse_seq.svh"
`include "sub_sequences/sync_pin/external_sync_pdcm_seq.svh"
`include "sub_sequences/sync_pin/measure_t_dsi3_sync_seq.svh"
`include "sub_sequences/sync_pin/mixed_external_internal_sync_seq.svh"
`include "sub_sequences/sync_pin/syncb_only_some_channels_seq.svh"
`include "sub_sequences/sync_pin/syncb_random_commands_seq.svh"
`include "sub_sequences/sync_pin/syncb_already_active_seq.svh"
`include "sub_sequences/sync_pin/syncb_during_running_crm_seq.svh"
`include "sub_sequences/sync_pin/syncb_sync_error_seq.svh"
`include "sub_sequences/sync_pin/syncb_short_pin_activation_seq.svh"

`include "sub_sequences/shift/apply_shift_while_in_pdcm_seq.svh"
`include "sub_sequences/shift/crm_shift_seq.svh"
`include "sub_sequences/shift/mix_starts_of_crm_seq.svh"
`include "sub_sequences/shift/pdcm_shift_seq.svh"
`include "sub_sequences/shift/pdcm_shift_sync_change_during_pdcm_seq.svh"
`include "sub_sequences/shift/pdcm_shift_sync_channel_1_before_0_seq.svh"
`include "sub_sequences/shift/pdcm_shift_sync_with_register_writes_seq.svh"
`include "sub_sequences/shift/pdcm_sync_change_while_pdcm_seq.svh"
`include "sub_sequences/shift/pdcm_sync_seq.svh"
`include "sub_sequences/shift/pdcm_sync_with_different_tdma_schemes_seq.svh"
`include "sub_sequences/shift/sync_between_pdcm_and_crm_seq.svh"
`include "sub_sequences/shift/discovery_mode_shift_seq.svh"

`include "sub_sequences/shut_off/dsi_enable_ignore_new_commands_seq.svh"
`include "sub_sequences/shut_off/dsi_enable_abort_crm_seq.sv"
`include "sub_sequences/shut_off/dsi_enable_abort_pdcm_seq.sv"
`include "sub_sequences/shut_off/dsi_enable_abort_command_queue_seq.svh"
`include "sub_sequences/shut_off/dsi_enable_abort_multi_packet_pdcm_seq.svh"
`include "sub_sequences/shut_off/dsi_enable_abort_discovery_mode_seq.svh"
`include "sub_sequences/shut_off/dsi_shut_off_and_check_crm_buffer_seq.svh"
`include "sub_sequences/shut_off/dsi_shut_off_and_check_pdcm_buffer_seq.svh"

`include "sub_sequences/tvl_base_shut_off_seq.svh"
`include "sub_sequences/overtemperature_shut_off_seq.svh"
`include "sub_sequences/overtemperature_status_seq.svh"
`include "sub_sequences/voltage_shut_off_seq.svh"
`include "sub_sequences/ldo_disable_shut_off_seq.svh"
`include "sub_sequences/tmr_out_seq.svh"
`include "sub_sequences/hardware_error_seq.svh"
`include "sub_sequences/sync_pin/sync_master_crm_seq.svh"
//
`include "ecc_error_base_seq.sv"
`include "sub_sequences/ecc/ecc_dsi3_receiver_rx_data_error_seq.svh"
`include "sub_sequences/ecc/ecc_dsi3_receiver_pdcm_to_ram_error_seq.svh"
`include "sub_sequences/ecc/ecc_dsi3_receiver_crm_to_ram_error_seq.svh"
`include "sub_sequences/ecc/ecc_dsi3_command_reading_error_seq.svh"
`include "sub_sequences/ecc/ecc_dsi3_crm_data_buffer_error_seq.svh"
`include "sub_sequences/ecc/ecc_dsi3_pdcm_data_buffer_error_seq.svh"
`include "sub_sequences/ecc/ecc_dsi3_command_buffer_error_seq.svh"
`include "sub_sequences/ecc/ecc_spi_command_buffer_error_seq.svh"
`include "sub_sequences/ecc/ecc_dsi3_tdma_error_seq.svh"
`include "sub_sequences/ecc/ecc_dsi3_transmit_data_error_seq.svh"
`include "sub_sequences/ecc/ecc_command_control_error_seq.svh"
`include "sub_sequences/ecc/ecc_spi_read_ram_data_error_seq.svh"
`include "sub_sequences/ecc/ecc_spi_read_dsi3_crm_data_error_seq.svh"
`include "sub_sequences/ecc/ecc_spi_read_dsi3_pdcm_data_error_seq.svh"
`include "sub_sequences/ecc/ecc_spi_received_data_error_seq.svh"
`include "sub_sequences/ecc/ecc_dsi3_data_high_low_error_seq.svh"
//`include "sub_sequences/ecc/ecc_dsi3_sync_error_seq.svh"

`include "sub_sequences/quiescent_current/quiescent_current_measurement_base_seq.svh"
`include "sub_sequences/quiescent_current/quiescent_current_seq.svh"
`include "sub_sequences/quiescent_current/manual_quiescent_current_measurement_seq.svh"

`include "applicative_pattern_seq.sv"
`include "applicative_pattern_ht_seq.sv"
`include "appl_examples_in_spec_seq.sv"
`include "debounce_times_seq.sv"
`include "dsi3_clear_command_buffer_seq.sv"
`include "dsi3_clear_data_buffer_seq.sv"
`include "dsi3_crm_seq.sv"
`include "dsi3_iload_seq.sv"
`include "dsi3_discovery_mode_seq.sv"
`include "dsi3_crm_ecc_1_bit_error_seq.sv"
`include "dsi3_crm_ecc_2_bit_error_seq.sv"
`include "dsi3_crm_timing_seq.sv"
`include "upload_tdma_seq.sv"
`include "dsi3_pdcm_seq.sv"
`include "dsi3_crc_seq.sv"
`include "dsi3_pdcm_timing_seq.sv"
`include "dsi3_sync_channels_seq.sv"
`include "dsi3_sync_pin_seq.sv"
`include "dsi3_sync_shift_seq.svh"
`include "dsi3_wait_seq.sv"
`include "jtag_test_seq.sv"
`include "register_access_seq.sv"
`include "shut_off_seq.svh"
`include "spi_errors_seq.svh"
`include "spi_framing_seq.svh"
`include "sub_sequences/base_irq_check_seq.sv"
`include "sub_sequences/interrupts/hierachical_irq_check_seq.sv"
`include "sub_sequences/interrupts/spi_base_irq_seq.sv"
`include "sub_sequences/interrupts/buf_base_irq_seq.sv"
`include "sub_sequences/interrupts/dsi_base_irq_seq.sv"
`include "sub_sequences/interrupts/buf_dsi_cmd_fe_irq_seq.sv"
`include "sub_sequences/interrupts/buf_dsi_crm_data_fe_irq_seq.sv"
`include "sub_sequences/interrupts/buf_dsi_pdcm_fe_irq_seq.sv"
`include "sub_sequences/interrupts/buf_spi_cmd_fe_irq_seq.sv"
`include "sub_sequences/interrupts/clkref_irq_seq.sv"
`include "sub_sequences/interrupts/dsi_com_err_irq_seq.sv"
`include "sub_sequences/interrupts/dsi_dmof_irq_seq.sv"
`include "sub_sequences/interrupts/dsi_dsiov_irq_seq.sv"
`include "sub_sequences/interrupts/dsi_dsiuv_irq_seq.sv"
`include "sub_sequences/interrupts/dsi_hw_fail_irq_seq.sv"
`include "sub_sequences/interrupts/dsi_iq_err_irq_seq.sv"
`include "sub_sequences/interrupts/dsi_sync_err_irq_seq.sv"
`include "sub_sequences/interrupts/hw_fail_irq_seq.sv"
`include "sub_sequences/interrupts/opt_fail_irq_seq.sv"
`include "sub_sequences/interrupts/reset_irq_seq.sv"
`include "sub_sequences/interrupts/spi_ali_err_irq_seq.sv"
`include "sub_sequences/interrupts/spi_cmd_ign_irq_seq.sv"
`include "sub_sequences/interrupts/spi_cmd_inc_irq_seq.sv"
`include "sub_sequences/interrupts/spi_crc_err_irq_seq.sv"
`include "sub_sequences/interrupts/spi_hw_fail_irq_seq.sv"
`include "sub_sequences/interrupts/supply_base_irq_seq.sv"
`include "sub_sequences/interrupts/supply_ldouv_irq_seq.sv"
`include "sub_sequences/interrupts/supply_ote_irq_seq.sv"
`include "sub_sequences/interrupts/supply_otw_irq_seq.sv"
`include "sub_sequences/interrupts/supply_ref_fail_irq_seq.sv"
`include "sub_sequences/interrupts/supply_vccuv_irq_seq.sv"
`include "interrupts_seq.sv"
`include "ic_startup_seq.sv"
`include "sram_bist_seq.sv"
`include "ic_status_word_seq.sv"
`include "uvm_register_sequences_seq.sv"
`include "otp_test_seq.sv"
`include "otp_trimming_seq.sv"
`include "otp_random_seq.sv"
`include "otp_pulse_width_seq.sv"
`include "ring_buffer_status_seq.sv"
`include "p52143_289_seq.sv"
`include "p52143_399_seq.sv"
`include "p52143_489_seq.sv"
`include "p52143_701_seq.sv"
`include "p52144_215_seq.sv"
//`include "pattern_compare_seq.sv"

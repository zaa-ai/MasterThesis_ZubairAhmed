/* ###   interface instances   ###################################################### */

Interrupt_Registers_IRQ_STAT_if Interrupt_Registers_IRQ_STAT (); 
Interrupt_Registers_IRQ_MASK_if Interrupt_Registers_IRQ_MASK (); 
Interrupt_Registers_ECC_IRQ_STAT_if Interrupt_Registers_ECC_IRQ_STAT (); 
Interrupt_Registers_ECC_IRQ_MASK_if Interrupt_Registers_ECC_IRQ_MASK (); 
Interrupt_Registers_ECC_CORR_IRQ_STAT_if Interrupt_Registers_ECC_CORR_IRQ_STAT (); 
Interrupt_Registers_ECC_CORR_IRQ_MASK_if Interrupt_Registers_ECC_CORR_IRQ_MASK (); 


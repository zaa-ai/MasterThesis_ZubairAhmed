
slave_timing[2][0].info_corner          = 0;
slave_timing[2][0].info_temp__j__       = 25;
slave_timing[2][0].info_i__quite_rec__  = 0.006000000;
slave_timing[2][0].info_dtr__ib__       = -1;
slave_timing[2][0].info_i__offset_rec__ = -0.001000000;
slave_timing[2][0].info_i__max_slave__  = 0.021000000;
slave_timing[2][0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][0].info_r__dsi_bus__    = 5.000;

slave_timing[2][0].t_rxd1[0][1] = 2835ns;
slave_timing[2][0].t_rxd1[1][0] = 2033ns;
slave_timing[2][0].t_rxd1[0][2] = 1958ns;
slave_timing[2][0].t_rxd1[2][0] = 2596ns;
slave_timing[2][0].t_rxd2[0][2] = 3161ns;
slave_timing[2][0].t_rxd2[2][0] = 1594ns;
slave_timing[2][0].t_rxd2[1][2] = 2856ns;
slave_timing[2][0].t_rxd2[2][1] = 2035ns;

slave_timing[2][1].info_corner          = 0;
slave_timing[2][1].info_temp__j__       = 25;
slave_timing[2][1].info_i__quite_rec__  = 0.006000000;
slave_timing[2][1].info_dtr__ib__       = -1;
slave_timing[2][1].info_i__offset_rec__ = 0.001000000;
slave_timing[2][1].info_i__max_slave__  = 0.021000000;
slave_timing[2][1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][1].info_r__dsi_bus__    = 5.000;

slave_timing[2][1].t_rxd1[0][1] = 2380ns;
slave_timing[2][1].t_rxd1[1][0] = 2410ns;
slave_timing[2][1].t_rxd1[0][2] = 1771ns;
slave_timing[2][1].t_rxd1[2][0] = 2835ns;
slave_timing[2][1].t_rxd2[0][2] = 2816ns;
slave_timing[2][1].t_rxd2[2][0] = 1803ns;
slave_timing[2][1].t_rxd2[1][2] = 2395ns;
slave_timing[2][1].t_rxd2[2][1] = 2418ns;

slave_timing[2][2].info_corner          = 0;
slave_timing[2][2].info_temp__j__       = 25;
slave_timing[2][2].info_i__quite_rec__  = 0.006000000;
slave_timing[2][2].info_dtr__ib__       = -1;
slave_timing[2][2].info_i__offset_rec__ = -0.001000000;
slave_timing[2][2].info_i__max_slave__  = 0.027000000;
slave_timing[2][2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][2].info_r__dsi_bus__    = 5.000;

slave_timing[2][2].t_rxd1[0][1] = 2398ns;
slave_timing[2][2].t_rxd1[1][0] = 2261ns;
slave_timing[2][2].t_rxd1[0][2] = 1781ns;
slave_timing[2][2].t_rxd1[2][0] = 2739ns;
slave_timing[2][2].t_rxd2[0][2] = 2548ns;
slave_timing[2][2].t_rxd2[2][0] = 1943ns;
slave_timing[2][2].t_rxd2[1][2] = 1982ns;
slave_timing[2][2].t_rxd2[2][1] = 2755ns;

slave_timing[2][3].info_corner          = 0;
slave_timing[2][3].info_temp__j__       = 25;
slave_timing[2][3].info_i__quite_rec__  = 0.006000000;
slave_timing[2][3].info_dtr__ib__       = -1;
slave_timing[2][3].info_i__offset_rec__ = 0.001000000;
slave_timing[2][3].info_i__max_slave__  = 0.027000000;
slave_timing[2][3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][3].info_r__dsi_bus__    = 5.000;

slave_timing[2][3].t_rxd1[0][1] = 2139ns;
slave_timing[2][3].t_rxd1[1][0] = 2537ns;
slave_timing[2][3].t_rxd1[0][2] = 1622ns;
slave_timing[2][3].t_rxd1[2][0] = 2933ns;
slave_timing[2][3].t_rxd2[0][2] = 2387ns;
slave_timing[2][3].t_rxd2[2][0] = 2069ns;
slave_timing[2][3].t_rxd2[1][2] = 1723ns;
slave_timing[2][3].t_rxd2[2][1] = 3244ns;

slave_timing[2][4].info_corner          = 0;
slave_timing[2][4].info_temp__j__       = 25;
slave_timing[2][4].info_i__quite_rec__  = 0.006000000;
slave_timing[2][4].info_dtr__ib__       = 1;
slave_timing[2][4].info_i__offset_rec__ = -0.001000000;
slave_timing[2][4].info_i__max_slave__  = 0.021000000;
slave_timing[2][4].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][4].info_r__dsi_bus__    = 5.000;

slave_timing[2][4].t_rxd1[0][1] = 2967ns;
slave_timing[2][4].t_rxd1[1][0] = 1979ns;
slave_timing[2][4].t_rxd1[0][2] = 1997ns;
slave_timing[2][4].t_rxd1[2][0] = 2560ns;
slave_timing[2][4].t_rxd2[0][2] = 3531ns;
slave_timing[2][4].t_rxd2[2][0] = 1479ns;
slave_timing[2][4].t_rxd2[1][2] = 3291ns;
slave_timing[2][4].t_rxd2[2][1] = 1866ns;

slave_timing[2][5].info_corner          = 0;
slave_timing[2][5].info_temp__j__       = 25;
slave_timing[2][5].info_i__quite_rec__  = 0.006000000;
slave_timing[2][5].info_dtr__ib__       = 1;
slave_timing[2][5].info_i__offset_rec__ = 0.001000000;
slave_timing[2][5].info_i__max_slave__  = 0.021000000;
slave_timing[2][5].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][5].info_r__dsi_bus__    = 5.000;

slave_timing[2][5].t_rxd1[0][1] = 2467ns;
slave_timing[2][5].t_rxd1[1][0] = 2350ns;
slave_timing[2][5].t_rxd1[0][2] = 1810ns;
slave_timing[2][5].t_rxd1[2][0] = 2800ns;
slave_timing[2][5].t_rxd2[0][2] = 2999ns;
slave_timing[2][5].t_rxd2[2][0] = 1705ns;
slave_timing[2][5].t_rxd2[1][2] = 2639ns;
slave_timing[2][5].t_rxd2[2][1] = 2225ns;

slave_timing[2][6].info_corner          = 0;
slave_timing[2][6].info_temp__j__       = 25;
slave_timing[2][6].info_i__quite_rec__  = 0.006000000;
slave_timing[2][6].info_dtr__ib__       = 1;
slave_timing[2][6].info_i__offset_rec__ = -0.001000000;
slave_timing[2][6].info_i__max_slave__  = 0.027000000;
slave_timing[2][6].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][6].info_r__dsi_bus__    = 5.000;

slave_timing[2][6].t_rxd1[0][1] = 2466ns;
slave_timing[2][6].t_rxd1[1][0] = 2221ns;
slave_timing[2][6].t_rxd1[0][2] = 1809ns;
slave_timing[2][6].t_rxd1[2][0] = 2712ns;
slave_timing[2][6].t_rxd2[0][2] = 2649ns;
slave_timing[2][6].t_rxd2[2][0] = 1874ns;
slave_timing[2][6].t_rxd2[1][2] = 2148ns;
slave_timing[2][6].t_rxd2[2][1] = 2579ns;

slave_timing[2][7].info_corner          = 0;
slave_timing[2][7].info_temp__j__       = 25;
slave_timing[2][7].info_i__quite_rec__  = 0.006000000;
slave_timing[2][7].info_dtr__ib__       = 1;
slave_timing[2][7].info_i__offset_rec__ = 0.001000000;
slave_timing[2][7].info_i__max_slave__  = 0.027000000;
slave_timing[2][7].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][7].info_r__dsi_bus__    = 5.000;

slave_timing[2][7].t_rxd1[0][1] = 2204ns;
slave_timing[2][7].t_rxd1[1][0] = 2490ns;
slave_timing[2][7].t_rxd1[0][2] = 1659ns;
slave_timing[2][7].t_rxd1[2][0] = 2899ns;
slave_timing[2][7].t_rxd2[0][2] = 2479ns;
slave_timing[2][7].t_rxd2[2][0] = 2000ns;
slave_timing[2][7].t_rxd2[1][2] = 1903ns;
slave_timing[2][7].t_rxd2[2][1] = 2931ns;

slave_timing[2][8].info_corner          = 0;
slave_timing[2][8].info_temp__j__       = 25;
slave_timing[2][8].info_i__quite_rec__  = 0.006000000;
slave_timing[2][8].info_dtr__ib__       = -1;
slave_timing[2][8].info_i__offset_rec__ = -0.001000000;
slave_timing[2][8].info_i__max_slave__  = 0.021000000;
slave_timing[2][8].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][8].info_r__dsi_bus__    = 5.000;

slave_timing[2][8].t_rxd1[0][1] = 3087ns;
slave_timing[2][8].t_rxd1[1][0] = 2240ns;
slave_timing[2][8].t_rxd1[0][2] = 2159ns;
slave_timing[2][8].t_rxd1[2][0] = 2828ns;
slave_timing[2][8].t_rxd2[0][2] = 3445ns;
slave_timing[2][8].t_rxd2[2][0] = 1780ns;
slave_timing[2][8].t_rxd2[1][2] = 3113ns;
slave_timing[2][8].t_rxd2[2][1] = 2244ns;

slave_timing[2][9].info_corner          = 0;
slave_timing[2][9].info_temp__j__       = 25;
slave_timing[2][9].info_i__quite_rec__  = 0.006000000;
slave_timing[2][9].info_dtr__ib__       = -1;
slave_timing[2][9].info_i__offset_rec__ = 0.001000000;
slave_timing[2][9].info_i__max_slave__  = 0.021000000;
slave_timing[2][9].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][9].info_r__dsi_bus__    = 5.000;

slave_timing[2][9].t_rxd1[0][1] = 2602ns;
slave_timing[2][9].t_rxd1[1][0] = 2632ns;
slave_timing[2][9].t_rxd1[0][2] = 1962ns;
slave_timing[2][9].t_rxd1[2][0] = 3089ns;
slave_timing[2][9].t_rxd2[0][2] = 3069ns;
slave_timing[2][9].t_rxd2[2][0] = 1993ns;
slave_timing[2][9].t_rxd2[1][2] = 2622ns;
slave_timing[2][9].t_rxd2[2][1] = 2638ns;

slave_timing[2][10].info_corner          = 0;
slave_timing[2][10].info_temp__j__       = 25;
slave_timing[2][10].info_i__quite_rec__  = 0.006000000;
slave_timing[2][10].info_dtr__ib__       = -1;
slave_timing[2][10].info_i__offset_rec__ = -0.001000000;
slave_timing[2][10].info_i__max_slave__  = 0.027000000;
slave_timing[2][10].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][10].info_r__dsi_bus__    = 5.000;

slave_timing[2][10].t_rxd1[0][1] = 2625ns;
slave_timing[2][10].t_rxd1[1][0] = 2486ns;
slave_timing[2][10].t_rxd1[0][2] = 1969ns;
slave_timing[2][10].t_rxd1[2][0] = 2984ns;
slave_timing[2][10].t_rxd2[0][2] = 2780ns;
slave_timing[2][10].t_rxd2[2][0] = 2141ns;
slave_timing[2][10].t_rxd2[1][2] = 2185ns;
slave_timing[2][10].t_rxd2[2][1] = 3005ns;

slave_timing[2][11].info_corner          = 0;
slave_timing[2][11].info_temp__j__       = 25;
slave_timing[2][11].info_i__quite_rec__  = 0.006000000;
slave_timing[2][11].info_dtr__ib__       = -1;
slave_timing[2][11].info_i__offset_rec__ = 0.001000000;
slave_timing[2][11].info_i__max_slave__  = 0.027000000;
slave_timing[2][11].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][11].info_r__dsi_bus__    = 5.000;

slave_timing[2][11].t_rxd1[0][1] = 2316ns;
slave_timing[2][11].t_rxd1[1][0] = 2803ns;
slave_timing[2][11].t_rxd1[0][2] = 1806ns;
slave_timing[2][11].t_rxd1[2][0] = 3224ns;
slave_timing[2][11].t_rxd2[0][2] = 2610ns;
slave_timing[2][11].t_rxd2[2][0] = 2290ns;
slave_timing[2][11].t_rxd2[1][2] = 1878ns;
slave_timing[2][11].t_rxd2[2][1] = 3646ns;

slave_timing[2][12].info_corner          = 0;
slave_timing[2][12].info_temp__j__       = 25;
slave_timing[2][12].info_i__quite_rec__  = 0.006000000;
slave_timing[2][12].info_dtr__ib__       = 1;
slave_timing[2][12].info_i__offset_rec__ = -0.001000000;
slave_timing[2][12].info_i__max_slave__  = 0.021000000;
slave_timing[2][12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][12].info_r__dsi_bus__    = 5.000;

slave_timing[2][12].t_rxd1[0][1] = 3237ns;
slave_timing[2][12].t_rxd1[1][0] = 2185ns;
slave_timing[2][12].t_rxd1[0][2] = 2202ns;
slave_timing[2][12].t_rxd1[2][0] = 2797ns;
slave_timing[2][12].t_rxd2[0][2] = 3857ns;
slave_timing[2][12].t_rxd2[2][0] = 1654ns;
slave_timing[2][12].t_rxd2[1][2] = 3585ns;
slave_timing[2][12].t_rxd2[2][1] = 2062ns;

slave_timing[2][13].info_corner          = 0;
slave_timing[2][13].info_temp__j__       = 25;
slave_timing[2][13].info_i__quite_rec__  = 0.006000000;
slave_timing[2][13].info_dtr__ib__       = 1;
slave_timing[2][13].info_i__offset_rec__ = 0.001000000;
slave_timing[2][13].info_i__max_slave__  = 0.021000000;
slave_timing[2][13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][13].info_r__dsi_bus__    = 5.000;

slave_timing[2][13].t_rxd1[0][1] = 2702ns;
slave_timing[2][13].t_rxd1[1][0] = 2566ns;
slave_timing[2][13].t_rxd1[0][2] = 2000ns;
slave_timing[2][13].t_rxd1[2][0] = 3053ns;
slave_timing[2][13].t_rxd2[0][2] = 3263ns;
slave_timing[2][13].t_rxd2[2][0] = 1893ns;
slave_timing[2][13].t_rxd2[1][2] = 2878ns;
slave_timing[2][13].t_rxd2[2][1] = 2452ns;

slave_timing[2][14].info_corner          = 0;
slave_timing[2][14].info_temp__j__       = 25;
slave_timing[2][14].info_i__quite_rec__  = 0.006000000;
slave_timing[2][14].info_dtr__ib__       = 1;
slave_timing[2][14].info_i__offset_rec__ = -0.001000000;
slave_timing[2][14].info_i__max_slave__  = 0.027000000;
slave_timing[2][14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][14].info_r__dsi_bus__    = 5.000;

slave_timing[2][14].t_rxd1[0][1] = 2700ns;
slave_timing[2][14].t_rxd1[1][0] = 2436ns;
slave_timing[2][14].t_rxd1[0][2] = 2006ns;
slave_timing[2][14].t_rxd1[2][0] = 2955ns;
slave_timing[2][14].t_rxd2[0][2] = 2889ns;
slave_timing[2][14].t_rxd2[2][0] = 2069ns;
slave_timing[2][14].t_rxd2[1][2] = 2361ns;
slave_timing[2][14].t_rxd2[2][1] = 2813ns;

slave_timing[2][15].info_corner          = 0;
slave_timing[2][15].info_temp__j__       = 25;
slave_timing[2][15].info_i__quite_rec__  = 0.006000000;
slave_timing[2][15].info_dtr__ib__       = 1;
slave_timing[2][15].info_i__offset_rec__ = 0.001000000;
slave_timing[2][15].info_i__max_slave__  = 0.027000000;
slave_timing[2][15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][15].info_r__dsi_bus__    = 5.000;

slave_timing[2][15].t_rxd1[0][1] = 2416ns;
slave_timing[2][15].t_rxd1[1][0] = 2715ns;
slave_timing[2][15].t_rxd1[0][2] = 1845ns;
slave_timing[2][15].t_rxd1[2][0] = 3155ns;
slave_timing[2][15].t_rxd2[0][2] = 2709ns;
slave_timing[2][15].t_rxd2[2][0] = 2202ns;
slave_timing[2][15].t_rxd2[1][2] = 2087ns;
slave_timing[2][15].t_rxd2[2][1] = 3198ns;

slave_timing[2][16].info_corner          = 0;
slave_timing[2][16].info_temp__j__       = 25;
slave_timing[2][16].info_i__quite_rec__  = 0.003000000;
slave_timing[2][16].info_dtr__ib__       = -1;
slave_timing[2][16].info_i__offset_rec__ = -0.001000000;
slave_timing[2][16].info_i__max_slave__  = 0.021000000;
slave_timing[2][16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][16].info_r__dsi_bus__    = 5.000;

slave_timing[2][16].t_rxd1[0][1] = 2809ns;
slave_timing[2][16].t_rxd1[1][0] = 2047ns;
slave_timing[2][16].t_rxd1[0][2] = 1951ns;
slave_timing[2][16].t_rxd1[2][0] = 2601ns;
slave_timing[2][16].t_rxd2[0][2] = 3148ns;
slave_timing[2][16].t_rxd2[2][0] = 1597ns;
slave_timing[2][16].t_rxd2[1][2] = 2832ns;
slave_timing[2][16].t_rxd2[2][1] = 2059ns;

slave_timing[2][17].info_corner          = 0;
slave_timing[2][17].info_temp__j__       = 25;
slave_timing[2][17].info_i__quite_rec__  = 0.003000000;
slave_timing[2][17].info_dtr__ib__       = -1;
slave_timing[2][17].info_i__offset_rec__ = 0.001000000;
slave_timing[2][17].info_i__max_slave__  = 0.021000000;
slave_timing[2][17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][17].info_r__dsi_bus__    = 5.000;

slave_timing[2][17].t_rxd1[0][1] = 2357ns;
slave_timing[2][17].t_rxd1[1][0] = 2420ns;
slave_timing[2][17].t_rxd1[0][2] = 1767ns;
slave_timing[2][17].t_rxd1[2][0] = 2850ns;
slave_timing[2][17].t_rxd2[0][2] = 2808ns;
slave_timing[2][17].t_rxd2[2][0] = 1809ns;
slave_timing[2][17].t_rxd2[1][2] = 2376ns;
slave_timing[2][17].t_rxd2[2][1] = 2427ns;

slave_timing[2][18].info_corner          = 0;
slave_timing[2][18].info_temp__j__       = 25;
slave_timing[2][18].info_i__quite_rec__  = 0.003000000;
slave_timing[2][18].info_dtr__ib__       = -1;
slave_timing[2][18].info_i__offset_rec__ = -0.001000000;
slave_timing[2][18].info_i__max_slave__  = 0.027000000;
slave_timing[2][18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][18].info_r__dsi_bus__    = 5.000;

slave_timing[2][18].t_rxd1[0][1] = 2382ns;
slave_timing[2][18].t_rxd1[1][0] = 2271ns;
slave_timing[2][18].t_rxd1[0][2] = 1787ns;
slave_timing[2][18].t_rxd1[2][0] = 2723ns;
slave_timing[2][18].t_rxd2[0][2] = 2555ns;
slave_timing[2][18].t_rxd2[2][0] = 1934ns;
slave_timing[2][18].t_rxd2[1][2] = 1967ns;
slave_timing[2][18].t_rxd2[2][1] = 2770ns;

slave_timing[2][19].info_corner          = 0;
slave_timing[2][19].info_temp__j__       = 25;
slave_timing[2][19].info_i__quite_rec__  = 0.003000000;
slave_timing[2][19].info_dtr__ib__       = -1;
slave_timing[2][19].info_i__offset_rec__ = 0.001000000;
slave_timing[2][19].info_i__max_slave__  = 0.027000000;
slave_timing[2][19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][19].info_r__dsi_bus__    = 5.000;

slave_timing[2][19].t_rxd1[0][1] = 2091ns;
slave_timing[2][19].t_rxd1[1][0] = 2582ns;
slave_timing[2][19].t_rxd1[0][2] = 1618ns;
slave_timing[2][19].t_rxd1[2][0] = 2966ns;
slave_timing[2][19].t_rxd2[0][2] = 2382ns;
slave_timing[2][19].t_rxd2[2][0] = 2083ns;
slave_timing[2][19].t_rxd2[1][2] = 1678ns;
slave_timing[2][19].t_rxd2[2][1] = 3375ns;

slave_timing[2][20].info_corner          = 0;
slave_timing[2][20].info_temp__j__       = 25;
slave_timing[2][20].info_i__quite_rec__  = 0.003000000;
slave_timing[2][20].info_dtr__ib__       = 1;
slave_timing[2][20].info_i__offset_rec__ = -0.001000000;
slave_timing[2][20].info_i__max_slave__  = 0.021000000;
slave_timing[2][20].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][20].info_r__dsi_bus__    = 5.000;

slave_timing[2][20].t_rxd1[0][1] = 2951ns;
slave_timing[2][20].t_rxd1[1][0] = 1992ns;
slave_timing[2][20].t_rxd1[0][2] = 1991ns;
slave_timing[2][20].t_rxd1[2][0] = 2565ns;
slave_timing[2][20].t_rxd2[0][2] = 3497ns;
slave_timing[2][20].t_rxd2[2][0] = 1479ns;
slave_timing[2][20].t_rxd2[1][2] = 3252ns;
slave_timing[2][20].t_rxd2[2][1] = 1879ns;

slave_timing[2][21].info_corner          = 0;
slave_timing[2][21].info_temp__j__       = 25;
slave_timing[2][21].info_i__quite_rec__  = 0.003000000;
slave_timing[2][21].info_dtr__ib__       = 1;
slave_timing[2][21].info_i__offset_rec__ = 0.001000000;
slave_timing[2][21].info_i__max_slave__  = 0.021000000;
slave_timing[2][21].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][21].info_r__dsi_bus__    = 5.000;

slave_timing[2][21].t_rxd1[0][1] = 2446ns;
slave_timing[2][21].t_rxd1[1][0] = 2367ns;
slave_timing[2][21].t_rxd1[0][2] = 1809ns;
slave_timing[2][21].t_rxd1[2][0] = 2810ns;
slave_timing[2][21].t_rxd2[0][2] = 2988ns;
slave_timing[2][21].t_rxd2[2][0] = 1713ns;
slave_timing[2][21].t_rxd2[1][2] = 2627ns;
slave_timing[2][21].t_rxd2[2][1] = 2239ns;

slave_timing[2][22].info_corner          = 0;
slave_timing[2][22].info_temp__j__       = 25;
slave_timing[2][22].info_i__quite_rec__  = 0.003000000;
slave_timing[2][22].info_dtr__ib__       = 1;
slave_timing[2][22].info_i__offset_rec__ = -0.001000000;
slave_timing[2][22].info_i__max_slave__  = 0.027000000;
slave_timing[2][22].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][22].info_r__dsi_bus__    = 5.000;

slave_timing[2][22].t_rxd1[0][1] = 2455ns;
slave_timing[2][22].t_rxd1[1][0] = 2230ns;
slave_timing[2][22].t_rxd1[0][2] = 1811ns;
slave_timing[2][22].t_rxd1[2][0] = 2716ns;
slave_timing[2][22].t_rxd2[0][2] = 2643ns;
slave_timing[2][22].t_rxd2[2][0] = 1880ns;
slave_timing[2][22].t_rxd2[1][2] = 2129ns;
slave_timing[2][22].t_rxd2[2][1] = 2591ns;

slave_timing[2][23].info_corner          = 0;
slave_timing[2][23].info_temp__j__       = 25;
slave_timing[2][23].info_i__quite_rec__  = 0.003000000;
slave_timing[2][23].info_dtr__ib__       = 1;
slave_timing[2][23].info_i__offset_rec__ = 0.001000000;
slave_timing[2][23].info_i__max_slave__  = 0.027000000;
slave_timing[2][23].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][23].info_r__dsi_bus__    = 5.000;

slave_timing[2][23].t_rxd1[0][1] = 2189ns;
slave_timing[2][23].t_rxd1[1][0] = 2495ns;
slave_timing[2][23].t_rxd1[0][2] = 1674ns;
slave_timing[2][23].t_rxd1[2][0] = 2904ns;
slave_timing[2][23].t_rxd2[0][2] = 2491ns;
slave_timing[2][23].t_rxd2[2][0] = 2005ns;
slave_timing[2][23].t_rxd2[1][2] = 1882ns;
slave_timing[2][23].t_rxd2[2][1] = 2944ns;

slave_timing[2][24].info_corner          = 0;
slave_timing[2][24].info_temp__j__       = 25;
slave_timing[2][24].info_i__quite_rec__  = 0.003000000;
slave_timing[2][24].info_dtr__ib__       = -1;
slave_timing[2][24].info_i__offset_rec__ = -0.001000000;
slave_timing[2][24].info_i__max_slave__  = 0.021000000;
slave_timing[2][24].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][24].info_r__dsi_bus__    = 5.000;

slave_timing[2][24].t_rxd1[0][1] = 3063ns;
slave_timing[2][24].t_rxd1[1][0] = 2259ns;
slave_timing[2][24].t_rxd1[0][2] = 2151ns;
slave_timing[2][24].t_rxd1[2][0] = 2838ns;
slave_timing[2][24].t_rxd2[0][2] = 3424ns;
slave_timing[2][24].t_rxd2[2][0] = 1782ns;
slave_timing[2][24].t_rxd2[1][2] = 3090ns;
slave_timing[2][24].t_rxd2[2][1] = 2260ns;

slave_timing[2][25].info_corner          = 0;
slave_timing[2][25].info_temp__j__       = 25;
slave_timing[2][25].info_i__quite_rec__  = 0.003000000;
slave_timing[2][25].info_dtr__ib__       = -1;
slave_timing[2][25].info_i__offset_rec__ = 0.001000000;
slave_timing[2][25].info_i__max_slave__  = 0.021000000;
slave_timing[2][25].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][25].info_r__dsi_bus__    = 5.000;

slave_timing[2][25].t_rxd1[0][1] = 2581ns;
slave_timing[2][25].t_rxd1[1][0] = 2647ns;
slave_timing[2][25].t_rxd1[0][2] = 1956ns;
slave_timing[2][25].t_rxd1[2][0] = 3100ns;
slave_timing[2][25].t_rxd2[0][2] = 3062ns;
slave_timing[2][25].t_rxd2[2][0] = 2001ns;
slave_timing[2][25].t_rxd2[1][2] = 2604ns;
slave_timing[2][25].t_rxd2[2][1] = 2649ns;

slave_timing[2][26].info_corner          = 0;
slave_timing[2][26].info_temp__j__       = 25;
slave_timing[2][26].info_i__quite_rec__  = 0.003000000;
slave_timing[2][26].info_dtr__ib__       = -1;
slave_timing[2][26].info_i__offset_rec__ = -0.001000000;
slave_timing[2][26].info_i__max_slave__  = 0.027000000;
slave_timing[2][26].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][26].info_r__dsi_bus__    = 5.000;

slave_timing[2][26].t_rxd1[0][1] = 2616ns;
slave_timing[2][26].t_rxd1[1][0] = 2487ns;
slave_timing[2][26].t_rxd1[0][2] = 1980ns;
slave_timing[2][26].t_rxd1[2][0] = 2969ns;
slave_timing[2][26].t_rxd2[0][2] = 2792ns;
slave_timing[2][26].t_rxd2[2][0] = 2133ns;
slave_timing[2][26].t_rxd2[1][2] = 2171ns;
slave_timing[2][26].t_rxd2[2][1] = 3015ns;

slave_timing[2][27].info_corner          = 0;
slave_timing[2][27].info_temp__j__       = 25;
slave_timing[2][27].info_i__quite_rec__  = 0.003000000;
slave_timing[2][27].info_dtr__ib__       = -1;
slave_timing[2][27].info_i__offset_rec__ = 0.001000000;
slave_timing[2][27].info_i__max_slave__  = 0.027000000;
slave_timing[2][27].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][27].info_r__dsi_bus__    = 5.000;

slave_timing[2][27].t_rxd1[0][1] = 2302ns;
slave_timing[2][27].t_rxd1[1][0] = 2819ns;
slave_timing[2][27].t_rxd1[0][2] = 1797ns;
slave_timing[2][27].t_rxd1[2][0] = 3225ns;
slave_timing[2][27].t_rxd2[0][2] = 2605ns;
slave_timing[2][27].t_rxd2[2][0] = 2291ns;
slave_timing[2][27].t_rxd2[1][2] = 1864ns;
slave_timing[2][27].t_rxd2[2][1] = 3581ns;

slave_timing[2][28].info_corner          = 0;
slave_timing[2][28].info_temp__j__       = 25;
slave_timing[2][28].info_i__quite_rec__  = 0.003000000;
slave_timing[2][28].info_dtr__ib__       = 1;
slave_timing[2][28].info_i__offset_rec__ = -0.001000000;
slave_timing[2][28].info_i__max_slave__  = 0.021000000;
slave_timing[2][28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][28].info_r__dsi_bus__    = 5.000;

slave_timing[2][28].t_rxd1[0][1] = 3198ns;
slave_timing[2][28].t_rxd1[1][0] = 2200ns;
slave_timing[2][28].t_rxd1[0][2] = 2196ns;
slave_timing[2][28].t_rxd1[2][0] = 2801ns;
slave_timing[2][28].t_rxd2[0][2] = 3821ns;
slave_timing[2][28].t_rxd2[2][0] = 1669ns;
slave_timing[2][28].t_rxd2[1][2] = 3533ns;
slave_timing[2][28].t_rxd2[2][1] = 2073ns;

slave_timing[2][29].info_corner          = 0;
slave_timing[2][29].info_temp__j__       = 25;
slave_timing[2][29].info_i__quite_rec__  = 0.003000000;
slave_timing[2][29].info_dtr__ib__       = 1;
slave_timing[2][29].info_i__offset_rec__ = 0.001000000;
slave_timing[2][29].info_i__max_slave__  = 0.021000000;
slave_timing[2][29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][29].info_r__dsi_bus__    = 5.000;

slave_timing[2][29].t_rxd1[0][1] = 2680ns;
slave_timing[2][29].t_rxd1[1][0] = 2577ns;
slave_timing[2][29].t_rxd1[0][2] = 2001ns;
slave_timing[2][29].t_rxd1[2][0] = 3057ns;
slave_timing[2][29].t_rxd2[0][2] = 3252ns;
slave_timing[2][29].t_rxd2[2][0] = 1891ns;
slave_timing[2][29].t_rxd2[1][2] = 2856ns;
slave_timing[2][29].t_rxd2[2][1] = 2452ns;

slave_timing[2][30].info_corner          = 0;
slave_timing[2][30].info_temp__j__       = 25;
slave_timing[2][30].info_i__quite_rec__  = 0.003000000;
slave_timing[2][30].info_dtr__ib__       = 1;
slave_timing[2][30].info_i__offset_rec__ = -0.001000000;
slave_timing[2][30].info_i__max_slave__  = 0.027000000;
slave_timing[2][30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][30].info_r__dsi_bus__    = 5.000;

slave_timing[2][30].t_rxd1[0][1] = 2682ns;
slave_timing[2][30].t_rxd1[1][0] = 2446ns;
slave_timing[2][30].t_rxd1[0][2] = 2003ns;
slave_timing[2][30].t_rxd1[2][0] = 2958ns;
slave_timing[2][30].t_rxd2[0][2] = 2881ns;
slave_timing[2][30].t_rxd2[2][0] = 2075ns;
slave_timing[2][30].t_rxd2[1][2] = 2343ns;
slave_timing[2][30].t_rxd2[2][1] = 2822ns;

slave_timing[2][31].info_corner          = 0;
slave_timing[2][31].info_temp__j__       = 25;
slave_timing[2][31].info_i__quite_rec__  = 0.003000000;
slave_timing[2][31].info_dtr__ib__       = 1;
slave_timing[2][31].info_i__offset_rec__ = 0.001000000;
slave_timing[2][31].info_i__max_slave__  = 0.027000000;
slave_timing[2][31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][31].info_r__dsi_bus__    = 5.000;

slave_timing[2][31].t_rxd1[0][1] = 2399ns;
slave_timing[2][31].t_rxd1[1][0] = 2727ns;
slave_timing[2][31].t_rxd1[0][2] = 1858ns;
slave_timing[2][31].t_rxd1[2][0] = 3165ns;
slave_timing[2][31].t_rxd2[0][2] = 2718ns;
slave_timing[2][31].t_rxd2[2][0] = 2209ns;
slave_timing[2][31].t_rxd2[1][2] = 2084ns;
slave_timing[2][31].t_rxd2[2][1] = 3207ns;

slave_timing[2][32].info_corner          = 0;
slave_timing[2][32].info_temp__j__       = 25;
slave_timing[2][32].info_i__quite_rec__  = 0.000000000;
slave_timing[2][32].info_dtr__ib__       = -1;
slave_timing[2][32].info_i__offset_rec__ = -0.001000000;
slave_timing[2][32].info_i__max_slave__  = 0.021000000;
slave_timing[2][32].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][32].info_r__dsi_bus__    = 5.000;

slave_timing[2][32].t_rxd1[0][1] = 2838ns;
slave_timing[2][32].t_rxd1[1][0] = 2029ns;
slave_timing[2][32].t_rxd1[0][2] = 1961ns;
slave_timing[2][32].t_rxd1[2][0] = 2594ns;
slave_timing[2][32].t_rxd2[0][2] = 3173ns;
slave_timing[2][32].t_rxd2[2][0] = 1594ns;
slave_timing[2][32].t_rxd2[1][2] = 2865ns;
slave_timing[2][32].t_rxd2[2][1] = 2033ns;

slave_timing[2][33].info_corner          = 0;
slave_timing[2][33].info_temp__j__       = 25;
slave_timing[2][33].info_i__quite_rec__  = 0.000000000;
slave_timing[2][33].info_dtr__ib__       = -1;
slave_timing[2][33].info_i__offset_rec__ = 0.001000000;
slave_timing[2][33].info_i__max_slave__  = 0.021000000;
slave_timing[2][33].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][33].info_r__dsi_bus__    = 5.000;

slave_timing[2][33].t_rxd1[0][1] = 2383ns;
slave_timing[2][33].t_rxd1[1][0] = 2407ns;
slave_timing[2][33].t_rxd1[0][2] = 1764ns;
slave_timing[2][33].t_rxd1[2][0] = 2836ns;
slave_timing[2][33].t_rxd2[0][2] = 2821ns;
slave_timing[2][33].t_rxd2[2][0] = 1800ns;
slave_timing[2][33].t_rxd2[1][2] = 2399ns;
slave_timing[2][33].t_rxd2[2][1] = 2413ns;

slave_timing[2][34].info_corner          = 0;
slave_timing[2][34].info_temp__j__       = 25;
slave_timing[2][34].info_i__quite_rec__  = 0.000000000;
slave_timing[2][34].info_dtr__ib__       = -1;
slave_timing[2][34].info_i__offset_rec__ = -0.001000000;
slave_timing[2][34].info_i__max_slave__  = 0.027000000;
slave_timing[2][34].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][34].info_r__dsi_bus__    = 5.000;

slave_timing[2][34].t_rxd1[0][1] = 2397ns;
slave_timing[2][34].t_rxd1[1][0] = 2264ns;
slave_timing[2][34].t_rxd1[0][2] = 1796ns;
slave_timing[2][34].t_rxd1[2][0] = 2721ns;
slave_timing[2][34].t_rxd2[0][2] = 2568ns;
slave_timing[2][34].t_rxd2[2][0] = 1929ns;
slave_timing[2][34].t_rxd2[1][2] = 1980ns;
slave_timing[2][34].t_rxd2[2][1] = 2755ns;

slave_timing[2][35].info_corner          = 0;
slave_timing[2][35].info_temp__j__       = 25;
slave_timing[2][35].info_i__quite_rec__  = 0.000000000;
slave_timing[2][35].info_dtr__ib__       = -1;
slave_timing[2][35].info_i__offset_rec__ = 0.001000000;
slave_timing[2][35].info_i__max_slave__  = 0.027000000;
slave_timing[2][35].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][35].info_r__dsi_bus__    = 5.000;

slave_timing[2][35].t_rxd1[0][1] = 2111ns;
slave_timing[2][35].t_rxd1[1][0] = 2569ns;
slave_timing[2][35].t_rxd1[0][2] = 1624ns;
slave_timing[2][35].t_rxd1[2][0] = 2954ns;
slave_timing[2][35].t_rxd2[0][2] = 2391ns;
slave_timing[2][35].t_rxd2[2][0] = 2078ns;
slave_timing[2][35].t_rxd2[1][2] = 1684ns;
slave_timing[2][35].t_rxd2[2][1] = 3327ns;

slave_timing[2][36].info_corner          = 0;
slave_timing[2][36].info_temp__j__       = 25;
slave_timing[2][36].info_i__quite_rec__  = 0.000000000;
slave_timing[2][36].info_dtr__ib__       = 1;
slave_timing[2][36].info_i__offset_rec__ = -0.001000000;
slave_timing[2][36].info_i__max_slave__  = 0.021000000;
slave_timing[2][36].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][36].info_r__dsi_bus__    = 5.000;

slave_timing[2][36].t_rxd1[0][1] = 3069ns;
slave_timing[2][36].t_rxd1[1][0] = 1936ns;
slave_timing[2][36].t_rxd1[0][2] = 2022ns;
slave_timing[2][36].t_rxd1[2][0] = 2532ns;
slave_timing[2][36].t_rxd2[0][2] = 3675ns;
slave_timing[2][36].t_rxd2[2][0] = 1437ns;
slave_timing[2][36].t_rxd2[1][2] = 3449ns;
slave_timing[2][36].t_rxd2[2][1] = 1814ns;

slave_timing[2][37].info_corner          = 0;
slave_timing[2][37].info_temp__j__       = 25;
slave_timing[2][37].info_i__quite_rec__  = 0.000000000;
slave_timing[2][37].info_dtr__ib__       = 1;
slave_timing[2][37].info_i__offset_rec__ = 0.001000000;
slave_timing[2][37].info_i__max_slave__  = 0.021000000;
slave_timing[2][37].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][37].info_r__dsi_bus__    = 5.000;

slave_timing[2][37].t_rxd1[0][1] = 2522ns;
slave_timing[2][37].t_rxd1[1][0] = 2302ns;
slave_timing[2][37].t_rxd1[0][2] = 1836ns;
slave_timing[2][37].t_rxd1[2][0] = 2766ns;
slave_timing[2][37].t_rxd2[0][2] = 3043ns;
slave_timing[2][37].t_rxd2[2][0] = 1672ns;
slave_timing[2][37].t_rxd2[1][2] = 2702ns;
slave_timing[2][37].t_rxd2[2][1] = 2179ns;

slave_timing[2][38].info_corner          = 0;
slave_timing[2][38].info_temp__j__       = 25;
slave_timing[2][38].info_i__quite_rec__  = 0.000000000;
slave_timing[2][38].info_dtr__ib__       = 1;
slave_timing[2][38].info_i__offset_rec__ = -0.001000000;
slave_timing[2][38].info_i__max_slave__  = 0.027000000;
slave_timing[2][38].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][38].info_r__dsi_bus__    = 5.000;

slave_timing[2][38].t_rxd1[0][1] = 2470ns;
slave_timing[2][38].t_rxd1[1][0] = 2215ns;
slave_timing[2][38].t_rxd1[0][2] = 1833ns;
slave_timing[2][38].t_rxd1[2][0] = 2686ns;
slave_timing[2][38].t_rxd2[0][2] = 2668ns;
slave_timing[2][38].t_rxd2[2][0] = 1858ns;
slave_timing[2][38].t_rxd2[1][2] = 2154ns;
slave_timing[2][38].t_rxd2[2][1] = 2568ns;

slave_timing[2][39].info_corner          = 0;
slave_timing[2][39].info_temp__j__       = 25;
slave_timing[2][39].info_i__quite_rec__  = 0.000000000;
slave_timing[2][39].info_dtr__ib__       = 1;
slave_timing[2][39].info_i__offset_rec__ = 0.001000000;
slave_timing[2][39].info_i__max_slave__  = 0.027000000;
slave_timing[2][39].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][39].info_r__dsi_bus__    = 5.000;

slave_timing[2][39].t_rxd1[0][1] = 2180ns;
slave_timing[2][39].t_rxd1[1][0] = 2509ns;
slave_timing[2][39].t_rxd1[0][2] = 1663ns;
slave_timing[2][39].t_rxd1[2][0] = 2918ns;
slave_timing[2][39].t_rxd2[0][2] = 2484ns;
slave_timing[2][39].t_rxd2[2][0] = 2009ns;
slave_timing[2][39].t_rxd2[1][2] = 1869ns;
slave_timing[2][39].t_rxd2[2][1] = 2970ns;

slave_timing[2][40].info_corner          = 0;
slave_timing[2][40].info_temp__j__       = 25;
slave_timing[2][40].info_i__quite_rec__  = 0.000000000;
slave_timing[2][40].info_dtr__ib__       = -1;
slave_timing[2][40].info_i__offset_rec__ = -0.001000000;
slave_timing[2][40].info_i__max_slave__  = 0.021000000;
slave_timing[2][40].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][40].info_r__dsi_bus__    = 5.000;

slave_timing[2][40].t_rxd1[0][1] = 3153ns;
slave_timing[2][40].t_rxd1[1][0] = 2207ns;
slave_timing[2][40].t_rxd1[0][2] = 2174ns;
slave_timing[2][40].t_rxd1[2][0] = 2809ns;
slave_timing[2][40].t_rxd2[0][2] = 3499ns;
slave_timing[2][40].t_rxd2[2][0] = 1752ns;
slave_timing[2][40].t_rxd2[1][2] = 3181ns;
slave_timing[2][40].t_rxd2[2][1] = 2207ns;

slave_timing[2][41].info_corner          = 0;
slave_timing[2][41].info_temp__j__       = 25;
slave_timing[2][41].info_i__quite_rec__  = 0.000000000;
slave_timing[2][41].info_dtr__ib__       = -1;
slave_timing[2][41].info_i__offset_rec__ = 0.001000000;
slave_timing[2][41].info_i__max_slave__  = 0.021000000;
slave_timing[2][41].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][41].info_r__dsi_bus__    = 5.000;

slave_timing[2][41].t_rxd1[0][1] = 2647ns;
slave_timing[2][41].t_rxd1[1][0] = 2589ns;
slave_timing[2][41].t_rxd1[0][2] = 1985ns;
slave_timing[2][41].t_rxd1[2][0] = 3053ns;
slave_timing[2][41].t_rxd2[0][2] = 3106ns;
slave_timing[2][41].t_rxd2[2][0] = 1970ns;
slave_timing[2][41].t_rxd2[1][2] = 2663ns;
slave_timing[2][41].t_rxd2[2][1] = 2592ns;

slave_timing[2][42].info_corner          = 0;
slave_timing[2][42].info_temp__j__       = 25;
slave_timing[2][42].info_i__quite_rec__  = 0.000000000;
slave_timing[2][42].info_dtr__ib__       = -1;
slave_timing[2][42].info_i__offset_rec__ = -0.001000000;
slave_timing[2][42].info_i__max_slave__  = 0.027000000;
slave_timing[2][42].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][42].info_r__dsi_bus__    = 5.000;

slave_timing[2][42].t_rxd1[0][1] = 2658ns;
slave_timing[2][42].t_rxd1[1][0] = 2448ns;
slave_timing[2][42].t_rxd1[0][2] = 1988ns;
slave_timing[2][42].t_rxd1[2][0] = 2962ns;
slave_timing[2][42].t_rxd2[0][2] = 2801ns;
slave_timing[2][42].t_rxd2[2][0] = 2128ns;
slave_timing[2][42].t_rxd2[1][2] = 2221ns;
slave_timing[2][42].t_rxd2[2][1] = 2958ns;

slave_timing[2][43].info_corner          = 0;
slave_timing[2][43].info_temp__j__       = 25;
slave_timing[2][43].info_i__quite_rec__  = 0.000000000;
slave_timing[2][43].info_dtr__ib__       = -1;
slave_timing[2][43].info_i__offset_rec__ = 0.001000000;
slave_timing[2][43].info_i__max_slave__  = 0.027000000;
slave_timing[2][43].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][43].info_r__dsi_bus__    = 5.000;

slave_timing[2][43].t_rxd1[0][1] = 2350ns;
slave_timing[2][43].t_rxd1[1][0] = 2770ns;
slave_timing[2][43].t_rxd1[0][2] = 1826ns;
slave_timing[2][43].t_rxd1[2][0] = 3190ns;
slave_timing[2][43].t_rxd2[0][2] = 2633ns;
slave_timing[2][43].t_rxd2[2][0] = 2273ns;
slave_timing[2][43].t_rxd2[1][2] = 1919ns;
slave_timing[2][43].t_rxd2[2][1] = 3528ns;

slave_timing[2][44].info_corner          = 0;
slave_timing[2][44].info_temp__j__       = 25;
slave_timing[2][44].info_i__quite_rec__  = 0.000000000;
slave_timing[2][44].info_dtr__ib__       = 1;
slave_timing[2][44].info_i__offset_rec__ = -0.001000000;
slave_timing[2][44].info_i__max_slave__  = 0.021000000;
slave_timing[2][44].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][44].info_r__dsi_bus__    = 5.000;

slave_timing[2][44].t_rxd1[0][1] = 3252ns;
slave_timing[2][44].t_rxd1[1][0] = 2182ns;
slave_timing[2][44].t_rxd1[0][2] = 2226ns;
slave_timing[2][44].t_rxd1[2][0] = 2767ns;
slave_timing[2][44].t_rxd2[0][2] = 4011ns;
slave_timing[2][44].t_rxd2[2][0] = 1615ns;
slave_timing[2][44].t_rxd2[1][2] = 3614ns;
slave_timing[2][44].t_rxd2[2][1] = 2049ns;

slave_timing[2][45].info_corner          = 0;
slave_timing[2][45].info_temp__j__       = 25;
slave_timing[2][45].info_i__quite_rec__  = 0.000000000;
slave_timing[2][45].info_dtr__ib__       = 1;
slave_timing[2][45].info_i__offset_rec__ = 0.001000000;
slave_timing[2][45].info_i__max_slave__  = 0.021000000;
slave_timing[2][45].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][45].info_r__dsi_bus__    = 5.000;

slave_timing[2][45].t_rxd1[0][1] = 2708ns;
slave_timing[2][45].t_rxd1[1][0] = 2560ns;
slave_timing[2][45].t_rxd1[0][2] = 2015ns;
slave_timing[2][45].t_rxd1[2][0] = 3042ns;
slave_timing[2][45].t_rxd2[0][2] = 3272ns;
slave_timing[2][45].t_rxd2[2][0] = 1882ns;
slave_timing[2][45].t_rxd2[1][2] = 2889ns;
slave_timing[2][45].t_rxd2[2][1] = 2436ns;

slave_timing[2][46].info_corner          = 0;
slave_timing[2][46].info_temp__j__       = 25;
slave_timing[2][46].info_i__quite_rec__  = 0.000000000;
slave_timing[2][46].info_dtr__ib__       = 1;
slave_timing[2][46].info_i__offset_rec__ = -0.001000000;
slave_timing[2][46].info_i__max_slave__  = 0.027000000;
slave_timing[2][46].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][46].info_r__dsi_bus__    = 5.000;

slave_timing[2][46].t_rxd1[0][1] = 2709ns;
slave_timing[2][46].t_rxd1[1][0] = 2426ns;
slave_timing[2][46].t_rxd1[0][2] = 2026ns;
slave_timing[2][46].t_rxd1[2][0] = 2930ns;
slave_timing[2][46].t_rxd2[0][2] = 2916ns;
slave_timing[2][46].t_rxd2[2][0] = 2052ns;
slave_timing[2][46].t_rxd2[1][2] = 2362ns;
slave_timing[2][46].t_rxd2[2][1] = 2802ns;

slave_timing[2][47].info_corner          = 0;
slave_timing[2][47].info_temp__j__       = 25;
slave_timing[2][47].info_i__quite_rec__  = 0.000000000;
slave_timing[2][47].info_dtr__ib__       = 1;
slave_timing[2][47].info_i__offset_rec__ = 0.001000000;
slave_timing[2][47].info_i__max_slave__  = 0.027000000;
slave_timing[2][47].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][47].info_r__dsi_bus__    = 5.000;

slave_timing[2][47].t_rxd1[0][1] = 2390ns;
slave_timing[2][47].t_rxd1[1][0] = 2745ns;
slave_timing[2][47].t_rxd1[0][2] = 1849ns;
slave_timing[2][47].t_rxd1[2][0] = 3176ns;
slave_timing[2][47].t_rxd2[0][2] = 2714ns;
slave_timing[2][47].t_rxd2[2][0] = 2213ns;
slave_timing[2][47].t_rxd2[1][2] = 2072ns;
slave_timing[2][47].t_rxd2[2][1] = 3230ns;

slave_timing[2][48].info_corner          = 0;
slave_timing[2][48].info_temp__j__       = 25;
slave_timing[2][48].info_i__quite_rec__  = 0.040000000;
slave_timing[2][48].info_dtr__ib__       = -1;
slave_timing[2][48].info_i__offset_rec__ = -0.001000000;
slave_timing[2][48].info_i__max_slave__  = 0.021000000;
slave_timing[2][48].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][48].info_r__dsi_bus__    = 5.000;

slave_timing[2][48].t_rxd1[0][1] = 2669ns;
slave_timing[2][48].t_rxd1[1][0] = 2149ns;
slave_timing[2][48].t_rxd1[0][2] = 1899ns;
slave_timing[2][48].t_rxd1[2][0] = 2665ns;
slave_timing[2][48].t_rxd2[0][2] = 3038ns;
slave_timing[2][48].t_rxd2[2][0] = 1663ns;
slave_timing[2][48].t_rxd2[1][2] = 2700ns;
slave_timing[2][48].t_rxd2[2][1] = 2150ns;

slave_timing[2][49].info_corner          = 0;
slave_timing[2][49].info_temp__j__       = 25;
slave_timing[2][49].info_i__quite_rec__  = 0.040000000;
slave_timing[2][49].info_dtr__ib__       = -1;
slave_timing[2][49].info_i__offset_rec__ = 0.001000000;
slave_timing[2][49].info_i__max_slave__  = 0.021000000;
slave_timing[2][49].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][49].info_r__dsi_bus__    = 5.000;

slave_timing[2][49].t_rxd1[0][1] = 2256ns;
slave_timing[2][49].t_rxd1[1][0] = 2534ns;
slave_timing[2][49].t_rxd1[0][2] = 1711ns;
slave_timing[2][49].t_rxd1[2][0] = 2926ns;
slave_timing[2][49].t_rxd2[0][2] = 2733ns;
slave_timing[2][49].t_rxd2[2][0] = 1848ns;
slave_timing[2][49].t_rxd2[1][2] = 2278ns;
slave_timing[2][49].t_rxd2[2][1] = 2531ns;

slave_timing[2][50].info_corner          = 0;
slave_timing[2][50].info_temp__j__       = 25;
slave_timing[2][50].info_i__quite_rec__  = 0.040000000;
slave_timing[2][50].info_dtr__ib__       = -1;
slave_timing[2][50].info_i__offset_rec__ = -0.001000000;
slave_timing[2][50].info_i__max_slave__  = 0.027000000;
slave_timing[2][50].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][50].info_r__dsi_bus__    = 5.000;

slave_timing[2][50].t_rxd1[0][1] = 2359ns;
slave_timing[2][50].t_rxd1[1][0] = 2306ns;
slave_timing[2][50].t_rxd1[0][2] = 1764ns;
slave_timing[2][50].t_rxd1[2][0] = 2761ns;
slave_timing[2][50].t_rxd2[0][2] = 2528ns;
slave_timing[2][50].t_rxd2[2][0] = 1957ns;
slave_timing[2][50].t_rxd2[1][2] = 1944ns;
slave_timing[2][50].t_rxd2[2][1] = 2790ns;

slave_timing[2][51].info_corner          = 0;
slave_timing[2][51].info_temp__j__       = 25;
slave_timing[2][51].info_i__quite_rec__  = 0.040000000;
slave_timing[2][51].info_dtr__ib__       = -1;
slave_timing[2][51].info_i__offset_rec__ = 0.001000000;
slave_timing[2][51].info_i__max_slave__  = 0.027000000;
slave_timing[2][51].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][51].info_r__dsi_bus__    = 5.000;

slave_timing[2][51].t_rxd1[0][1] = 2107ns;
slave_timing[2][51].t_rxd1[1][0] = 2581ns;
slave_timing[2][51].t_rxd1[0][2] = 1618ns;
slave_timing[2][51].t_rxd1[2][0] = 2963ns;
slave_timing[2][51].t_rxd2[0][2] = 2387ns;
slave_timing[2][51].t_rxd2[2][0] = 2080ns;
slave_timing[2][51].t_rxd2[1][2] = 1688ns;
slave_timing[2][51].t_rxd2[2][1] = 3345ns;

slave_timing[2][52].info_corner          = 0;
slave_timing[2][52].info_temp__j__       = 25;
slave_timing[2][52].info_i__quite_rec__  = 0.040000000;
slave_timing[2][52].info_dtr__ib__       = 1;
slave_timing[2][52].info_i__offset_rec__ = -0.001000000;
slave_timing[2][52].info_i__max_slave__  = 0.021000000;
slave_timing[2][52].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][52].info_r__dsi_bus__    = 5.000;

slave_timing[2][52].t_rxd1[0][1] = 3011ns;
slave_timing[2][52].t_rxd1[1][0] = 1957ns;
slave_timing[2][52].t_rxd1[0][2] = 2008ns;
slave_timing[2][52].t_rxd1[2][0] = 2548ns;
slave_timing[2][52].t_rxd2[0][2] = 3585ns;
slave_timing[2][52].t_rxd2[2][0] = 1455ns;
slave_timing[2][52].t_rxd2[1][2] = 3350ns;
slave_timing[2][52].t_rxd2[2][1] = 1842ns;

slave_timing[2][53].info_corner          = 0;
slave_timing[2][53].info_temp__j__       = 25;
slave_timing[2][53].info_i__quite_rec__  = 0.040000000;
slave_timing[2][53].info_dtr__ib__       = 1;
slave_timing[2][53].info_i__offset_rec__ = 0.001000000;
slave_timing[2][53].info_i__max_slave__  = 0.021000000;
slave_timing[2][53].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][53].info_r__dsi_bus__    = 5.000;

slave_timing[2][53].t_rxd1[0][1] = 2491ns;
slave_timing[2][53].t_rxd1[1][0] = 2326ns;
slave_timing[2][53].t_rxd1[0][2] = 1824ns;
slave_timing[2][53].t_rxd1[2][0] = 2783ns;
slave_timing[2][53].t_rxd2[0][2] = 3013ns;
slave_timing[2][53].t_rxd2[2][0] = 1690ns;
slave_timing[2][53].t_rxd2[1][2] = 2652ns;
slave_timing[2][53].t_rxd2[2][1] = 2213ns;

slave_timing[2][54].info_corner          = 0;
slave_timing[2][54].info_temp__j__       = 25;
slave_timing[2][54].info_i__quite_rec__  = 0.040000000;
slave_timing[2][54].info_dtr__ib__       = 1;
slave_timing[2][54].info_i__offset_rec__ = -0.001000000;
slave_timing[2][54].info_i__max_slave__  = 0.027000000;
slave_timing[2][54].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][54].info_r__dsi_bus__    = 5.000;

slave_timing[2][54].t_rxd1[0][1] = 2526ns;
slave_timing[2][54].t_rxd1[1][0] = 2174ns;
slave_timing[2][54].t_rxd1[0][2] = 1836ns;
slave_timing[2][54].t_rxd1[2][0] = 2680ns;
slave_timing[2][54].t_rxd2[0][2] = 2678ns;
slave_timing[2][54].t_rxd2[2][0] = 1852ns;
slave_timing[2][54].t_rxd2[1][2] = 2191ns;
slave_timing[2][54].t_rxd2[2][1] = 2526ns;

slave_timing[2][55].info_corner          = 0;
slave_timing[2][55].info_temp__j__       = 25;
slave_timing[2][55].info_i__quite_rec__  = 0.040000000;
slave_timing[2][55].info_dtr__ib__       = 1;
slave_timing[2][55].info_i__offset_rec__ = 0.001000000;
slave_timing[2][55].info_i__max_slave__  = 0.027000000;
slave_timing[2][55].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][55].info_r__dsi_bus__    = 5.000;

slave_timing[2][55].t_rxd1[0][1] = 2213ns;
slave_timing[2][55].t_rxd1[1][0] = 2473ns;
slave_timing[2][55].t_rxd1[0][2] = 1685ns;
slave_timing[2][55].t_rxd1[2][0] = 2883ns;
slave_timing[2][55].t_rxd2[0][2] = 2499ns;
slave_timing[2][55].t_rxd2[2][0] = 1991ns;
slave_timing[2][55].t_rxd2[1][2] = 1909ns;
slave_timing[2][55].t_rxd2[2][1] = 2901ns;

slave_timing[2][56].info_corner          = 0;
slave_timing[2][56].info_temp__j__       = 25;
slave_timing[2][56].info_i__quite_rec__  = 0.040000000;
slave_timing[2][56].info_dtr__ib__       = -1;
slave_timing[2][56].info_i__offset_rec__ = -0.001000000;
slave_timing[2][56].info_i__max_slave__  = 0.021000000;
slave_timing[2][56].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][56].info_r__dsi_bus__    = 5.000;

slave_timing[2][56].t_rxd1[0][1] = 2913ns;
slave_timing[2][56].t_rxd1[1][0] = 2364ns;
slave_timing[2][56].t_rxd1[0][2] = 2101ns;
slave_timing[2][56].t_rxd1[2][0] = 2903ns;
slave_timing[2][56].t_rxd2[0][2] = 3308ns;
slave_timing[2][56].t_rxd2[2][0] = 1846ns;
slave_timing[2][56].t_rxd2[1][2] = 2935ns;
slave_timing[2][56].t_rxd2[2][1] = 2362ns;

slave_timing[2][57].info_corner          = 0;
slave_timing[2][57].info_temp__j__       = 25;
slave_timing[2][57].info_i__quite_rec__  = 0.040000000;
slave_timing[2][57].info_dtr__ib__       = -1;
slave_timing[2][57].info_i__offset_rec__ = 0.001000000;
slave_timing[2][57].info_i__max_slave__  = 0.021000000;
slave_timing[2][57].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][57].info_r__dsi_bus__    = 5.000;

slave_timing[2][57].t_rxd1[0][1] = 2477ns;
slave_timing[2][57].t_rxd1[1][0] = 2765ns;
slave_timing[2][57].t_rxd1[0][2] = 1902ns;
slave_timing[2][57].t_rxd1[2][0] = 3189ns;
slave_timing[2][57].t_rxd2[0][2] = 2990ns;
slave_timing[2][57].t_rxd2[2][0] = 2052ns;
slave_timing[2][57].t_rxd2[1][2] = 2493ns;
slave_timing[2][57].t_rxd2[2][1] = 2768ns;

slave_timing[2][58].info_corner          = 0;
slave_timing[2][58].info_temp__j__       = 25;
slave_timing[2][58].info_i__quite_rec__  = 0.040000000;
slave_timing[2][58].info_dtr__ib__       = -1;
slave_timing[2][58].info_i__offset_rec__ = -0.001000000;
slave_timing[2][58].info_i__max_slave__  = 0.027000000;
slave_timing[2][58].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][58].info_r__dsi_bus__    = 5.000;

slave_timing[2][58].t_rxd1[0][1] = 2582ns;
slave_timing[2][58].t_rxd1[1][0] = 2529ns;
slave_timing[2][58].t_rxd1[0][2] = 1954ns;
slave_timing[2][58].t_rxd1[2][0] = 3011ns;
slave_timing[2][58].t_rxd2[0][2] = 2762ns;
slave_timing[2][58].t_rxd2[2][0] = 2157ns;
slave_timing[2][58].t_rxd2[1][2] = 2150ns;
slave_timing[2][58].t_rxd2[2][1] = 3048ns;

slave_timing[2][59].info_corner          = 0;
slave_timing[2][59].info_temp__j__       = 25;
slave_timing[2][59].info_i__quite_rec__  = 0.040000000;
slave_timing[2][59].info_dtr__ib__       = -1;
slave_timing[2][59].info_i__offset_rec__ = 0.001000000;
slave_timing[2][59].info_i__max_slave__  = 0.027000000;
slave_timing[2][59].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][59].info_r__dsi_bus__    = 5.000;

slave_timing[2][59].t_rxd1[0][1] = 2310ns;
slave_timing[2][59].t_rxd1[1][0] = 2811ns;
slave_timing[2][59].t_rxd1[0][2] = 1802ns;
slave_timing[2][59].t_rxd1[2][0] = 3230ns;
slave_timing[2][59].t_rxd2[0][2] = 2612ns;
slave_timing[2][59].t_rxd2[2][0] = 2289ns;
slave_timing[2][59].t_rxd2[1][2] = 1873ns;
slave_timing[2][59].t_rxd2[2][1] = 3661ns;

slave_timing[2][60].info_corner          = 0;
slave_timing[2][60].info_temp__j__       = 25;
slave_timing[2][60].info_i__quite_rec__  = 0.040000000;
slave_timing[2][60].info_dtr__ib__       = 1;
slave_timing[2][60].info_i__offset_rec__ = -0.001000000;
slave_timing[2][60].info_i__max_slave__  = 0.021000000;
slave_timing[2][60].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][60].info_r__dsi_bus__    = 5.000;

slave_timing[2][60].t_rxd1[0][1] = 3270ns;
slave_timing[2][60].t_rxd1[1][0] = 2165ns;
slave_timing[2][60].t_rxd1[0][2] = 2212ns;
slave_timing[2][60].t_rxd1[2][0] = 2780ns;
slave_timing[2][60].t_rxd2[0][2] = 3911ns;
slave_timing[2][60].t_rxd2[2][0] = 1640ns;
slave_timing[2][60].t_rxd2[1][2] = 3648ns;
slave_timing[2][60].t_rxd2[2][1] = 2042ns;

slave_timing[2][61].info_corner          = 0;
slave_timing[2][61].info_temp__j__       = 25;
slave_timing[2][61].info_i__quite_rec__  = 0.040000000;
slave_timing[2][61].info_dtr__ib__       = 1;
slave_timing[2][61].info_i__offset_rec__ = 0.001000000;
slave_timing[2][61].info_i__max_slave__  = 0.021000000;
slave_timing[2][61].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][61].info_r__dsi_bus__    = 5.000;

slave_timing[2][61].t_rxd1[0][1] = 2722ns;
slave_timing[2][61].t_rxd1[1][0] = 2555ns;
slave_timing[2][61].t_rxd1[0][2] = 2023ns;
slave_timing[2][61].t_rxd1[2][0] = 3033ns;
slave_timing[2][61].t_rxd2[0][2] = 3285ns;
slave_timing[2][61].t_rxd2[2][0] = 1884ns;
slave_timing[2][61].t_rxd2[1][2] = 2904ns;
slave_timing[2][61].t_rxd2[2][1] = 2417ns;

slave_timing[2][62].info_corner          = 0;
slave_timing[2][62].info_temp__j__       = 25;
slave_timing[2][62].info_i__quite_rec__  = 0.040000000;
slave_timing[2][62].info_dtr__ib__       = 1;
slave_timing[2][62].info_i__offset_rec__ = -0.001000000;
slave_timing[2][62].info_i__max_slave__  = 0.027000000;
slave_timing[2][62].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][62].info_r__dsi_bus__    = 5.000;

slave_timing[2][62].t_rxd1[0][1] = 2716ns;
slave_timing[2][62].t_rxd1[1][0] = 2419ns;
slave_timing[2][62].t_rxd1[0][2] = 2017ns;
slave_timing[2][62].t_rxd1[2][0] = 2940ns;
slave_timing[2][62].t_rxd2[0][2] = 2899ns;
slave_timing[2][62].t_rxd2[2][0] = 2061ns;
slave_timing[2][62].t_rxd2[1][2] = 2371ns;
slave_timing[2][62].t_rxd2[2][1] = 2793ns;

slave_timing[2][63].info_corner          = 0;
slave_timing[2][63].info_temp__j__       = 25;
slave_timing[2][63].info_i__quite_rec__  = 0.040000000;
slave_timing[2][63].info_dtr__ib__       = 1;
slave_timing[2][63].info_i__offset_rec__ = 0.001000000;
slave_timing[2][63].info_i__max_slave__  = 0.027000000;
slave_timing[2][63].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][63].info_r__dsi_bus__    = 5.000;

slave_timing[2][63].t_rxd1[0][1] = 2434ns;
slave_timing[2][63].t_rxd1[1][0] = 2698ns;
slave_timing[2][63].t_rxd1[0][2] = 1873ns;
slave_timing[2][63].t_rxd1[2][0] = 3139ns;
slave_timing[2][63].t_rxd2[0][2] = 2736ns;
slave_timing[2][63].t_rxd2[2][0] = 2196ns;
slave_timing[2][63].t_rxd2[1][2] = 2109ns;
slave_timing[2][63].t_rxd2[2][1] = 3159ns;

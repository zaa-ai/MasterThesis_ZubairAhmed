
slave_timing[1][96+0].info_corner          = 4;
slave_timing[1][96+0].info_temp__j__       = 125;
slave_timing[1][96+0].info_i__quite_rec__  = 0.006000000;
slave_timing[1][96+0].info_dtr__ib__       = -1;
slave_timing[1][96+0].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+0].info_i__max_slave__  = 0.023000000;
slave_timing[1][96+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][96+0].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+0].t_rxd1[0][1] = 1657ns;
slave_timing[1][96+0].t_rxd1[1][0] = 1634ns;
slave_timing[1][96+0].t_rxd1[0][2] = 1245ns;
slave_timing[1][96+0].t_rxd1[2][0] = 1977ns;
slave_timing[1][96+0].t_rxd2[0][2] = 2012ns;
slave_timing[1][96+0].t_rxd2[2][0] = 1246ns;
slave_timing[1][96+0].t_rxd2[1][2] = 1696ns;
slave_timing[1][96+0].t_rxd2[2][1] = 1633ns;

slave_timing[1][96+1].info_corner          = 4;
slave_timing[1][96+1].info_temp__j__       = 125;
slave_timing[1][96+1].info_i__quite_rec__  = 0.006000000;
slave_timing[1][96+1].info_dtr__ib__       = -1;
slave_timing[1][96+1].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+1].info_i__max_slave__  = 0.025000000;
slave_timing[1][96+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][96+1].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+1].t_rxd1[0][1] = 1592ns;
slave_timing[1][96+1].t_rxd1[1][0] = 1682ns;
slave_timing[1][96+1].t_rxd1[0][2] = 1208ns;
slave_timing[1][96+1].t_rxd1[2][0] = 2010ns;
slave_timing[1][96+1].t_rxd2[0][2] = 1887ns;
slave_timing[1][96+1].t_rxd2[2][0] = 1329ns;
slave_timing[1][96+1].t_rxd2[1][2] = 1517ns;
slave_timing[1][96+1].t_rxd2[2][1] = 1799ns;

slave_timing[1][96+2].info_corner          = 4;
slave_timing[1][96+2].info_temp__j__       = 125;
slave_timing[1][96+2].info_i__quite_rec__  = 0.006000000;
slave_timing[1][96+2].info_dtr__ib__       = 1;
slave_timing[1][96+2].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+2].info_i__max_slave__  = 0.023000000;
slave_timing[1][96+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][96+2].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+2].t_rxd1[0][1] = 1667ns;
slave_timing[1][96+2].t_rxd1[1][0] = 1587ns;
slave_timing[1][96+2].t_rxd1[0][2] = 1244ns;
slave_timing[1][96+2].t_rxd1[2][0] = 1929ns;
slave_timing[1][96+2].t_rxd2[0][2] = 2083ns;
slave_timing[1][96+2].t_rxd2[2][0] = 1178ns;
slave_timing[1][96+2].t_rxd2[1][2] = 1805ns;
slave_timing[1][96+2].t_rxd2[2][1] = 1511ns;

slave_timing[1][96+3].info_corner          = 4;
slave_timing[1][96+3].info_temp__j__       = 125;
slave_timing[1][96+3].info_i__quite_rec__  = 0.006000000;
slave_timing[1][96+3].info_dtr__ib__       = 1;
slave_timing[1][96+3].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+3].info_i__max_slave__  = 0.025000000;
slave_timing[1][96+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][96+3].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+3].t_rxd1[0][1] = 1600ns;
slave_timing[1][96+3].t_rxd1[1][0] = 1634ns;
slave_timing[1][96+3].t_rxd1[0][2] = 1208ns;
slave_timing[1][96+3].t_rxd1[2][0] = 1962ns;
slave_timing[1][96+3].t_rxd2[0][2] = 1938ns;
slave_timing[1][96+3].t_rxd2[2][0] = 1267ns;
slave_timing[1][96+3].t_rxd2[1][2] = 1606ns;
slave_timing[1][96+3].t_rxd2[2][1] = 1678ns;

slave_timing[1][96+4].info_corner          = 4;
slave_timing[1][96+4].info_temp__j__       = 125;
slave_timing[1][96+4].info_i__quite_rec__  = 0.006000000;
slave_timing[1][96+4].info_dtr__ib__       = -1;
slave_timing[1][96+4].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+4].info_i__max_slave__  = 0.023000000;
slave_timing[1][96+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][96+4].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+4].t_rxd1[0][1] = 1840ns;
slave_timing[1][96+4].t_rxd1[1][0] = 1766ns;
slave_timing[1][96+4].t_rxd1[0][2] = 1389ns;
slave_timing[1][96+4].t_rxd1[2][0] = 2099ns;
slave_timing[1][96+4].t_rxd2[0][2] = 2055ns;
slave_timing[1][96+4].t_rxd2[2][0] = 1277ns;
slave_timing[1][96+4].t_rxd2[1][2] = 1714ns;
slave_timing[1][96+4].t_rxd2[2][1] = 1654ns;

slave_timing[1][96+5].info_corner          = 4;
slave_timing[1][96+5].info_temp__j__       = 125;
slave_timing[1][96+5].info_i__quite_rec__  = 0.006000000;
slave_timing[1][96+5].info_dtr__ib__       = -1;
slave_timing[1][96+5].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+5].info_i__max_slave__  = 0.025000000;
slave_timing[1][96+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][96+5].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+5].t_rxd1[0][1] = 1768ns;
slave_timing[1][96+5].t_rxd1[1][0] = 1813ns;
slave_timing[1][96+5].t_rxd1[0][2] = 1352ns;
slave_timing[1][96+5].t_rxd1[2][0] = 2130ns;
slave_timing[1][96+5].t_rxd2[0][2] = 1935ns;
slave_timing[1][96+5].t_rxd2[2][0] = 1358ns;
slave_timing[1][96+5].t_rxd2[1][2] = 1540ns;
slave_timing[1][96+5].t_rxd2[2][1] = 1818ns;

slave_timing[1][96+6].info_corner          = 4;
slave_timing[1][96+6].info_temp__j__       = 125;
slave_timing[1][96+6].info_i__quite_rec__  = 0.006000000;
slave_timing[1][96+6].info_dtr__ib__       = 1;
slave_timing[1][96+6].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+6].info_i__max_slave__  = 0.023000000;
slave_timing[1][96+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][96+6].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+6].t_rxd1[0][1] = 1847ns;
slave_timing[1][96+6].t_rxd1[1][0] = 1713ns;
slave_timing[1][96+6].t_rxd1[0][2] = 1383ns;
slave_timing[1][96+6].t_rxd1[2][0] = 2044ns;
slave_timing[1][96+6].t_rxd2[0][2] = 2119ns;
slave_timing[1][96+6].t_rxd2[2][0] = 1205ns;
slave_timing[1][96+6].t_rxd2[1][2] = 1822ns;
slave_timing[1][96+6].t_rxd2[2][1] = 1536ns;

slave_timing[1][96+7].info_corner          = 4;
slave_timing[1][96+7].info_temp__j__       = 125;
slave_timing[1][96+7].info_i__quite_rec__  = 0.006000000;
slave_timing[1][96+7].info_dtr__ib__       = 1;
slave_timing[1][96+7].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+7].info_i__max_slave__  = 0.025000000;
slave_timing[1][96+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][96+7].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+7].t_rxd1[0][1] = 1773ns;
slave_timing[1][96+7].t_rxd1[1][0] = 1759ns;
slave_timing[1][96+7].t_rxd1[0][2] = 1348ns;
slave_timing[1][96+7].t_rxd1[2][0] = 2076ns;
slave_timing[1][96+7].t_rxd2[0][2] = 1977ns;
slave_timing[1][96+7].t_rxd2[2][0] = 1295ns;
slave_timing[1][96+7].t_rxd2[1][2] = 1627ns;
slave_timing[1][96+7].t_rxd2[2][1] = 1678ns;

slave_timing[1][96+8].info_corner          = 4;
slave_timing[1][96+8].info_temp__j__       = 125;
slave_timing[1][96+8].info_i__quite_rec__  = 0.003000000;
slave_timing[1][96+8].info_dtr__ib__       = -1;
slave_timing[1][96+8].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+8].info_i__max_slave__  = 0.023000000;
slave_timing[1][96+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][96+8].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+8].t_rxd1[0][1] = 1621ns;
slave_timing[1][96+8].t_rxd1[1][0] = 1602ns;
slave_timing[1][96+8].t_rxd1[0][2] = 1220ns;
slave_timing[1][96+8].t_rxd1[2][0] = 1929ns;
slave_timing[1][96+8].t_rxd2[0][2] = 1971ns;
slave_timing[1][96+8].t_rxd2[2][0] = 1222ns;
slave_timing[1][96+8].t_rxd2[1][2] = 1669ns;
slave_timing[1][96+8].t_rxd2[2][1] = 1595ns;

slave_timing[1][96+9].info_corner          = 4;
slave_timing[1][96+9].info_temp__j__       = 125;
slave_timing[1][96+9].info_i__quite_rec__  = 0.003000000;
slave_timing[1][96+9].info_dtr__ib__       = -1;
slave_timing[1][96+9].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+9].info_i__max_slave__  = 0.025000000;
slave_timing[1][96+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][96+9].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+9].t_rxd1[0][1] = 1557ns;
slave_timing[1][96+9].t_rxd1[1][0] = 1646ns;
slave_timing[1][96+9].t_rxd1[0][2] = 1183ns;
slave_timing[1][96+9].t_rxd1[2][0] = 1960ns;
slave_timing[1][96+9].t_rxd2[0][2] = 1849ns;
slave_timing[1][96+9].t_rxd2[2][0] = 1303ns;
slave_timing[1][96+9].t_rxd2[1][2] = 1496ns;
slave_timing[1][96+9].t_rxd2[2][1] = 1758ns;

slave_timing[1][96+10].info_corner          = 4;
slave_timing[1][96+10].info_temp__j__       = 125;
slave_timing[1][96+10].info_i__quite_rec__  = 0.003000000;
slave_timing[1][96+10].info_dtr__ib__       = 1;
slave_timing[1][96+10].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+10].info_i__max_slave__  = 0.023000000;
slave_timing[1][96+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][96+10].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+10].t_rxd1[0][1] = 1644ns;
slave_timing[1][96+10].t_rxd1[1][0] = 1556ns;
slave_timing[1][96+10].t_rxd1[0][2] = 1225ns;
slave_timing[1][96+10].t_rxd1[2][0] = 1886ns;
slave_timing[1][96+10].t_rxd2[0][2] = 2038ns;
slave_timing[1][96+10].t_rxd2[2][0] = 1142ns;
slave_timing[1][96+10].t_rxd2[1][2] = 1775ns;
slave_timing[1][96+10].t_rxd2[2][1] = 1465ns;

slave_timing[1][96+11].info_corner          = 4;
slave_timing[1][96+11].info_temp__j__       = 125;
slave_timing[1][96+11].info_i__quite_rec__  = 0.003000000;
slave_timing[1][96+11].info_dtr__ib__       = 1;
slave_timing[1][96+11].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+11].info_i__max_slave__  = 0.025000000;
slave_timing[1][96+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][96+11].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+11].t_rxd1[0][1] = 1576ns;
slave_timing[1][96+11].t_rxd1[1][0] = 1606ns;
slave_timing[1][96+11].t_rxd1[0][2] = 1188ns;
slave_timing[1][96+11].t_rxd1[2][0] = 1917ns;
slave_timing[1][96+11].t_rxd2[0][2] = 1897ns;
slave_timing[1][96+11].t_rxd2[2][0] = 1232ns;
slave_timing[1][96+11].t_rxd2[1][2] = 1582ns;
slave_timing[1][96+11].t_rxd2[2][1] = 1626ns;

slave_timing[1][96+12].info_corner          = 4;
slave_timing[1][96+12].info_temp__j__       = 125;
slave_timing[1][96+12].info_i__quite_rec__  = 0.003000000;
slave_timing[1][96+12].info_dtr__ib__       = -1;
slave_timing[1][96+12].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+12].info_i__max_slave__  = 0.023000000;
slave_timing[1][96+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][96+12].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+12].t_rxd1[0][1] = 1821ns;
slave_timing[1][96+12].t_rxd1[1][0] = 1735ns;
slave_timing[1][96+12].t_rxd1[0][2] = 1374ns;
slave_timing[1][96+12].t_rxd1[2][0] = 2050ns;
slave_timing[1][96+12].t_rxd2[0][2] = 2006ns;
slave_timing[1][96+12].t_rxd2[2][0] = 1249ns;
slave_timing[1][96+12].t_rxd2[1][2] = 1687ns;
slave_timing[1][96+12].t_rxd2[2][1] = 1616ns;

slave_timing[1][96+13].info_corner          = 4;
slave_timing[1][96+13].info_temp__j__       = 125;
slave_timing[1][96+13].info_i__quite_rec__  = 0.003000000;
slave_timing[1][96+13].info_dtr__ib__       = -1;
slave_timing[1][96+13].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+13].info_i__max_slave__  = 0.025000000;
slave_timing[1][96+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][96+13].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+13].t_rxd1[0][1] = 1751ns;
slave_timing[1][96+13].t_rxd1[1][0] = 1778ns;
slave_timing[1][96+13].t_rxd1[0][2] = 1338ns;
slave_timing[1][96+13].t_rxd1[2][0] = 2081ns;
slave_timing[1][96+13].t_rxd2[0][2] = 1892ns;
slave_timing[1][96+13].t_rxd2[2][0] = 1331ns;
slave_timing[1][96+13].t_rxd2[1][2] = 1519ns;
slave_timing[1][96+13].t_rxd2[2][1] = 1777ns;

slave_timing[1][96+14].info_corner          = 4;
slave_timing[1][96+14].info_temp__j__       = 125;
slave_timing[1][96+14].info_i__quite_rec__  = 0.003000000;
slave_timing[1][96+14].info_dtr__ib__       = 1;
slave_timing[1][96+14].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+14].info_i__max_slave__  = 0.023000000;
slave_timing[1][96+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][96+14].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+14].t_rxd1[0][1] = 1838ns;
slave_timing[1][96+14].t_rxd1[1][0] = 1688ns;
slave_timing[1][96+14].t_rxd1[0][2] = 1380ns;
slave_timing[1][96+14].t_rxd1[2][0] = 2001ns;
slave_timing[1][96+14].t_rxd2[0][2] = 2069ns;
slave_timing[1][96+14].t_rxd2[2][0] = 1169ns;
slave_timing[1][96+14].t_rxd2[1][2] = 1792ns;
slave_timing[1][96+14].t_rxd2[2][1] = 1487ns;

slave_timing[1][96+15].info_corner          = 4;
slave_timing[1][96+15].info_temp__j__       = 125;
slave_timing[1][96+15].info_i__quite_rec__  = 0.003000000;
slave_timing[1][96+15].info_dtr__ib__       = 1;
slave_timing[1][96+15].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+15].info_i__max_slave__  = 0.025000000;
slave_timing[1][96+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][96+15].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+15].t_rxd1[0][1] = 1766ns;
slave_timing[1][96+15].t_rxd1[1][0] = 1734ns;
slave_timing[1][96+15].t_rxd1[0][2] = 1338ns;
slave_timing[1][96+15].t_rxd1[2][0] = 2030ns;
slave_timing[1][96+15].t_rxd2[0][2] = 1933ns;
slave_timing[1][96+15].t_rxd2[2][0] = 1259ns;
slave_timing[1][96+15].t_rxd2[1][2] = 1602ns;
slave_timing[1][96+15].t_rxd2[2][1] = 1646ns;

slave_timing[1][96+16].info_corner          = 4;
slave_timing[1][96+16].info_temp__j__       = 125;
slave_timing[1][96+16].info_i__quite_rec__  = 0.000000000;
slave_timing[1][96+16].info_dtr__ib__       = -1;
slave_timing[1][96+16].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+16].info_i__max_slave__  = 0.023000000;
slave_timing[1][96+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][96+16].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+16].t_rxd1[0][1] = 1599ns;
slave_timing[1][96+16].t_rxd1[1][0] = 1569ns;
slave_timing[1][96+16].t_rxd1[0][2] = 1203ns;
slave_timing[1][96+16].t_rxd1[2][0] = 1883ns;
slave_timing[1][96+16].t_rxd2[0][2] = 1923ns;
slave_timing[1][96+16].t_rxd2[2][0] = 1187ns;
slave_timing[1][96+16].t_rxd2[1][2] = 1634ns;
slave_timing[1][96+16].t_rxd2[2][1] = 1548ns;

slave_timing[1][96+17].info_corner          = 4;
slave_timing[1][96+17].info_temp__j__       = 125;
slave_timing[1][96+17].info_i__quite_rec__  = 0.000000000;
slave_timing[1][96+17].info_dtr__ib__       = -1;
slave_timing[1][96+17].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+17].info_i__max_slave__  = 0.025000000;
slave_timing[1][96+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][96+17].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+17].t_rxd1[0][1] = 1538ns;
slave_timing[1][96+17].t_rxd1[1][0] = 1615ns;
slave_timing[1][96+17].t_rxd1[0][2] = 1169ns;
slave_timing[1][96+17].t_rxd1[2][0] = 1912ns;
slave_timing[1][96+17].t_rxd2[0][2] = 1805ns;
slave_timing[1][96+17].t_rxd2[2][0] = 1268ns;
slave_timing[1][96+17].t_rxd2[1][2] = 1466ns;
slave_timing[1][96+17].t_rxd2[2][1] = 1703ns;

slave_timing[1][96+18].info_corner          = 4;
slave_timing[1][96+18].info_temp__j__       = 125;
slave_timing[1][96+18].info_i__quite_rec__  = 0.000000000;
slave_timing[1][96+18].info_dtr__ib__       = 1;
slave_timing[1][96+18].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+18].info_i__max_slave__  = 0.023000000;
slave_timing[1][96+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][96+18].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+18].t_rxd1[0][1] = 1615ns;
slave_timing[1][96+18].t_rxd1[1][0] = 1529ns;
slave_timing[1][96+18].t_rxd1[0][2] = 1204ns;
slave_timing[1][96+18].t_rxd1[2][0] = 1847ns;
slave_timing[1][96+18].t_rxd2[0][2] = 1993ns;
slave_timing[1][96+18].t_rxd2[2][0] = 1112ns;
slave_timing[1][96+18].t_rxd2[1][2] = 1740ns;
slave_timing[1][96+18].t_rxd2[2][1] = 1427ns;

slave_timing[1][96+19].info_corner          = 4;
slave_timing[1][96+19].info_temp__j__       = 125;
slave_timing[1][96+19].info_i__quite_rec__  = 0.000000000;
slave_timing[1][96+19].info_dtr__ib__       = 1;
slave_timing[1][96+19].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+19].info_i__max_slave__  = 0.025000000;
slave_timing[1][96+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][96+19].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+19].t_rxd1[0][1] = 1550ns;
slave_timing[1][96+19].t_rxd1[1][0] = 1572ns;
slave_timing[1][96+19].t_rxd1[0][2] = 1168ns;
slave_timing[1][96+19].t_rxd1[2][0] = 1878ns;
slave_timing[1][96+19].t_rxd2[0][2] = 1855ns;
slave_timing[1][96+19].t_rxd2[2][0] = 1200ns;
slave_timing[1][96+19].t_rxd2[1][2] = 1546ns;
slave_timing[1][96+19].t_rxd2[2][1] = 1583ns;

slave_timing[1][96+20].info_corner          = 4;
slave_timing[1][96+20].info_temp__j__       = 125;
slave_timing[1][96+20].info_i__quite_rec__  = 0.000000000;
slave_timing[1][96+20].info_dtr__ib__       = -1;
slave_timing[1][96+20].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+20].info_i__max_slave__  = 0.023000000;
slave_timing[1][96+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][96+20].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+20].t_rxd1[0][1] = 1821ns;
slave_timing[1][96+20].t_rxd1[1][0] = 1703ns;
slave_timing[1][96+20].t_rxd1[0][2] = 1377ns;
slave_timing[1][96+20].t_rxd1[2][0] = 1999ns;
slave_timing[1][96+20].t_rxd2[0][2] = 1956ns;
slave_timing[1][96+20].t_rxd2[2][0] = 1216ns;
slave_timing[1][96+20].t_rxd2[1][2] = 1653ns;
slave_timing[1][96+20].t_rxd2[2][1] = 1568ns;

slave_timing[1][96+21].info_corner          = 4;
slave_timing[1][96+21].info_temp__j__       = 125;
slave_timing[1][96+21].info_i__quite_rec__  = 0.000000000;
slave_timing[1][96+21].info_dtr__ib__       = -1;
slave_timing[1][96+21].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+21].info_i__max_slave__  = 0.025000000;
slave_timing[1][96+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][96+21].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+21].t_rxd1[0][1] = 1752ns;
slave_timing[1][96+21].t_rxd1[1][0] = 1745ns;
slave_timing[1][96+21].t_rxd1[0][2] = 1339ns;
slave_timing[1][96+21].t_rxd1[2][0] = 2027ns;
slave_timing[1][96+21].t_rxd2[0][2] = 1843ns;
slave_timing[1][96+21].t_rxd2[2][0] = 1294ns;
slave_timing[1][96+21].t_rxd2[1][2] = 1493ns;
slave_timing[1][96+21].t_rxd2[2][1] = 1701ns;

slave_timing[1][96+22].info_corner          = 4;
slave_timing[1][96+22].info_temp__j__       = 125;
slave_timing[1][96+22].info_i__quite_rec__  = 0.000000000;
slave_timing[1][96+22].info_dtr__ib__       = 1;
slave_timing[1][96+22].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+22].info_i__max_slave__  = 0.023000000;
slave_timing[1][96+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][96+22].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+22].t_rxd1[0][1] = 1833ns;
slave_timing[1][96+22].t_rxd1[1][0] = 1656ns;
slave_timing[1][96+22].t_rxd1[0][2] = 1376ns;
slave_timing[1][96+22].t_rxd1[2][0] = 1960ns;
slave_timing[1][96+22].t_rxd2[0][2] = 2017ns;
slave_timing[1][96+22].t_rxd2[2][0] = 1139ns;
slave_timing[1][96+22].t_rxd2[1][2] = 1754ns;
slave_timing[1][96+22].t_rxd2[2][1] = 1433ns;

slave_timing[1][96+23].info_corner          = 4;
slave_timing[1][96+23].info_temp__j__       = 125;
slave_timing[1][96+23].info_i__quite_rec__  = 0.000000000;
slave_timing[1][96+23].info_dtr__ib__       = 1;
slave_timing[1][96+23].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+23].info_i__max_slave__  = 0.025000000;
slave_timing[1][96+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][96+23].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+23].t_rxd1[0][1] = 1762ns;
slave_timing[1][96+23].t_rxd1[1][0] = 1698ns;
slave_timing[1][96+23].t_rxd1[0][2] = 1338ns;
slave_timing[1][96+23].t_rxd1[2][0] = 1990ns;
slave_timing[1][96+23].t_rxd2[0][2] = 1887ns;
slave_timing[1][96+23].t_rxd2[2][0] = 1228ns;
slave_timing[1][96+23].t_rxd2[1][2] = 1566ns;
slave_timing[1][96+23].t_rxd2[2][1] = 1585ns;

slave_timing[1][96+24].info_corner          = 4;
slave_timing[1][96+24].info_temp__j__       = 125;
slave_timing[1][96+24].info_i__quite_rec__  = 0.040000000;
slave_timing[1][96+24].info_dtr__ib__       = -1;
slave_timing[1][96+24].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+24].info_i__max_slave__  = 0.023000000;
slave_timing[1][96+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][96+24].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+24].t_rxd1[0][1] = 1725ns;
slave_timing[1][96+24].t_rxd1[1][0] = 1699ns;
slave_timing[1][96+24].t_rxd1[0][2] = 1331ns;
slave_timing[1][96+24].t_rxd1[2][0] = 2111ns;
slave_timing[1][96+24].t_rxd2[0][2] = 2302ns;
slave_timing[1][96+24].t_rxd2[2][0] = 1450ns;
slave_timing[1][96+24].t_rxd2[1][2] = 1955ns;
slave_timing[1][96+24].t_rxd2[2][1] = 1888ns;

slave_timing[1][96+25].info_corner          = 4;
slave_timing[1][96+25].info_temp__j__       = 125;
slave_timing[1][96+25].info_i__quite_rec__  = 0.040000000;
slave_timing[1][96+25].info_dtr__ib__       = -1;
slave_timing[1][96+25].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+25].info_i__max_slave__  = 0.025000000;
slave_timing[1][96+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][96+25].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+25].t_rxd1[0][1] = 1665ns;
slave_timing[1][96+25].t_rxd1[1][0] = 1756ns;
slave_timing[1][96+25].t_rxd1[0][2] = 1297ns;
slave_timing[1][96+25].t_rxd1[2][0] = 2154ns;
slave_timing[1][96+25].t_rxd2[0][2] = 2164ns;
slave_timing[1][96+25].t_rxd2[2][0] = 1538ns;
slave_timing[1][96+25].t_rxd2[1][2] = 1758ns;
slave_timing[1][96+25].t_rxd2[2][1] = 2076ns;

slave_timing[1][96+26].info_corner          = 4;
slave_timing[1][96+26].info_temp__j__       = 125;
slave_timing[1][96+26].info_i__quite_rec__  = 0.040000000;
slave_timing[1][96+26].info_dtr__ib__       = 1;
slave_timing[1][96+26].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+26].info_i__max_slave__  = 0.023000000;
slave_timing[1][96+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][96+26].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+26].t_rxd1[0][1] = 1775ns;
slave_timing[1][96+26].t_rxd1[1][0] = 1653ns;
slave_timing[1][96+26].t_rxd1[0][2] = 1357ns;
slave_timing[1][96+26].t_rxd1[2][0] = 2077ns;
slave_timing[1][96+26].t_rxd2[0][2] = 2419ns;
slave_timing[1][96+26].t_rxd2[2][0] = 1375ns;
slave_timing[1][96+26].t_rxd2[1][2] = 2107ns;
slave_timing[1][96+26].t_rxd2[2][1] = 1754ns;

slave_timing[1][96+27].info_corner          = 4;
slave_timing[1][96+27].info_temp__j__       = 125;
slave_timing[1][96+27].info_i__quite_rec__  = 0.040000000;
slave_timing[1][96+27].info_dtr__ib__       = 1;
slave_timing[1][96+27].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+27].info_i__max_slave__  = 0.025000000;
slave_timing[1][96+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][96+27].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+27].t_rxd1[0][1] = 1708ns;
slave_timing[1][96+27].t_rxd1[1][0] = 1711ns;
slave_timing[1][96+27].t_rxd1[0][2] = 1321ns;
slave_timing[1][96+27].t_rxd1[2][0] = 2118ns;
slave_timing[1][96+27].t_rxd2[0][2] = 2251ns;
slave_timing[1][96+27].t_rxd2[2][0] = 1470ns;
slave_timing[1][96+27].t_rxd2[1][2] = 1886ns;
slave_timing[1][96+27].t_rxd2[2][1] = 1938ns;

slave_timing[1][96+28].info_corner          = 4;
slave_timing[1][96+28].info_temp__j__       = 125;
slave_timing[1][96+28].info_i__quite_rec__  = 0.040000000;
slave_timing[1][96+28].info_dtr__ib__       = -1;
slave_timing[1][96+28].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+28].info_i__max_slave__  = 0.023000000;
slave_timing[1][96+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][96+28].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+28].t_rxd1[0][1] = 1820ns;
slave_timing[1][96+28].t_rxd1[1][0] = 2123ns;
slave_timing[1][96+28].t_rxd1[0][2] = 1445ns;
slave_timing[1][96+28].t_rxd1[2][0] = 2990ns;
slave_timing[1][96+28].t_rxd2[0][2] = 3228ns;
slave_timing[1][96+28].t_rxd2[2][0] = 1973ns;
slave_timing[1][96+28].t_rxd2[1][2] = 2769ns;
slave_timing[1][96+28].t_rxd2[2][1] = 2717ns;

slave_timing[1][96+29].info_corner          = 4;
slave_timing[1][96+29].info_temp__j__       = 125;
slave_timing[1][96+29].info_i__quite_rec__  = 0.040000000;
slave_timing[1][96+29].info_dtr__ib__       = -1;
slave_timing[1][96+29].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+29].info_i__max_slave__  = 0.025000000;
slave_timing[1][96+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][96+29].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+29].t_rxd1[0][1] = 1763ns;
slave_timing[1][96+29].t_rxd1[1][0] = 2223ns;
slave_timing[1][96+29].t_rxd1[0][2] = 1412ns;
slave_timing[1][96+29].t_rxd1[2][0] = 3094ns;
slave_timing[1][96+29].t_rxd2[0][2] = 2956ns;
slave_timing[1][96+29].t_rxd2[2][0] = 2114ns;
slave_timing[1][96+29].t_rxd2[1][2] = 2426ns;
slave_timing[1][96+29].t_rxd2[2][1] = 3116ns;

slave_timing[1][96+30].info_corner          = 4;
slave_timing[1][96+30].info_temp__j__       = 125;
slave_timing[1][96+30].info_i__quite_rec__  = 0.040000000;
slave_timing[1][96+30].info_dtr__ib__       = 1;
slave_timing[1][96+30].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+30].info_i__max_slave__  = 0.023000000;
slave_timing[1][96+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][96+30].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+30].t_rxd1[0][1] = 1863ns;
slave_timing[1][96+30].t_rxd1[1][0] = 2005ns;
slave_timing[1][96+30].t_rxd1[0][2] = 1468ns;
slave_timing[1][96+30].t_rxd1[2][0] = 2866ns;
slave_timing[1][96+30].t_rxd2[0][2] = 3471ns;
slave_timing[1][96+30].t_rxd2[2][0] = 1854ns;
slave_timing[1][96+30].t_rxd2[1][2] = 3058ns;
slave_timing[1][96+30].t_rxd2[2][1] = 2452ns;

slave_timing[1][96+31].info_corner          = 4;
slave_timing[1][96+31].info_temp__j__       = 125;
slave_timing[1][96+31].info_i__quite_rec__  = 0.040000000;
slave_timing[1][96+31].info_dtr__ib__       = 1;
slave_timing[1][96+31].info_i__offset_rec__ = 0.000000000;
slave_timing[1][96+31].info_i__max_slave__  = 0.025000000;
slave_timing[1][96+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][96+31].info_r__dsi_bus__    = 5.000;

slave_timing[1][96+31].t_rxd1[0][1] = 1800ns;
slave_timing[1][96+31].t_rxd1[1][0] = 2109ns;
slave_timing[1][96+31].t_rxd1[0][2] = 1432ns;
slave_timing[1][96+31].t_rxd1[2][0] = 2968ns;
slave_timing[1][96+31].t_rxd2[0][2] = 3116ns;
slave_timing[1][96+31].t_rxd2[2][0] = 2005ns;
slave_timing[1][96+31].t_rxd2[1][2] = 2642ns;
slave_timing[1][96+31].t_rxd2[2][1] = 2804ns;

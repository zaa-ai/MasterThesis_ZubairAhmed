
slave_timing[1][160+0].info_corner          = 2;
slave_timing[1][160+0].info_temp__j__       = -40;
slave_timing[1][160+0].info_i__quite_rec__  = 0.006000000;
slave_timing[1][160+0].info_dtr__ib__       = -1;
slave_timing[1][160+0].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+0].info_i__max_slave__  = 0.023000000;
slave_timing[1][160+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][160+0].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+0].t_rxd1[0][1] = 1657ns;
slave_timing[1][160+0].t_rxd1[1][0] = 1664ns;
slave_timing[1][160+0].t_rxd1[0][2] = 1246ns;
slave_timing[1][160+0].t_rxd1[2][0] = 2023ns;
slave_timing[1][160+0].t_rxd2[0][2] = 1997ns;
slave_timing[1][160+0].t_rxd2[2][0] = 1246ns;
slave_timing[1][160+0].t_rxd2[1][2] = 1639ns;
slave_timing[1][160+0].t_rxd2[2][1] = 1652ns;

slave_timing[1][160+1].info_corner          = 2;
slave_timing[1][160+1].info_temp__j__       = -40;
slave_timing[1][160+1].info_i__quite_rec__  = 0.006000000;
slave_timing[1][160+1].info_dtr__ib__       = -1;
slave_timing[1][160+1].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+1].info_i__max_slave__  = 0.025000000;
slave_timing[1][160+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][160+1].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+1].t_rxd1[0][1] = 1594ns;
slave_timing[1][160+1].t_rxd1[1][0] = 1715ns;
slave_timing[1][160+1].t_rxd1[0][2] = 1210ns;
slave_timing[1][160+1].t_rxd1[2][0] = 2057ns;
slave_timing[1][160+1].t_rxd2[0][2] = 1878ns;
slave_timing[1][160+1].t_rxd2[2][0] = 1329ns;
slave_timing[1][160+1].t_rxd2[1][2] = 1463ns;
slave_timing[1][160+1].t_rxd2[2][1] = 1825ns;

slave_timing[1][160+2].info_corner          = 2;
slave_timing[1][160+2].info_temp__j__       = -40;
slave_timing[1][160+2].info_i__quite_rec__  = 0.006000000;
slave_timing[1][160+2].info_dtr__ib__       = 1;
slave_timing[1][160+2].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+2].info_i__max_slave__  = 0.023000000;
slave_timing[1][160+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][160+2].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+2].t_rxd1[0][1] = 1705ns;
slave_timing[1][160+2].t_rxd1[1][0] = 1627ns;
slave_timing[1][160+2].t_rxd1[0][2] = 1271ns;
slave_timing[1][160+2].t_rxd1[2][0] = 1995ns;
slave_timing[1][160+2].t_rxd2[0][2] = 2107ns;
slave_timing[1][160+2].t_rxd2[2][0] = 1176ns;
slave_timing[1][160+2].t_rxd2[1][2] = 1787ns;
slave_timing[1][160+2].t_rxd2[2][1] = 1525ns;

slave_timing[1][160+3].info_corner          = 2;
slave_timing[1][160+3].info_temp__j__       = -40;
slave_timing[1][160+3].info_i__quite_rec__  = 0.006000000;
slave_timing[1][160+3].info_dtr__ib__       = 1;
slave_timing[1][160+3].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+3].info_i__max_slave__  = 0.025000000;
slave_timing[1][160+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][160+3].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+3].t_rxd1[0][1] = 1636ns;
slave_timing[1][160+3].t_rxd1[1][0] = 1677ns;
slave_timing[1][160+3].t_rxd1[0][2] = 1235ns;
slave_timing[1][160+3].t_rxd1[2][0] = 2031ns;
slave_timing[1][160+3].t_rxd2[0][2] = 1962ns;
slave_timing[1][160+3].t_rxd2[2][0] = 1267ns;
slave_timing[1][160+3].t_rxd2[1][2] = 1590ns;
slave_timing[1][160+3].t_rxd2[2][1] = 1695ns;

slave_timing[1][160+4].info_corner          = 2;
slave_timing[1][160+4].info_temp__j__       = -40;
slave_timing[1][160+4].info_i__quite_rec__  = 0.006000000;
slave_timing[1][160+4].info_dtr__ib__       = -1;
slave_timing[1][160+4].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+4].info_i__max_slave__  = 0.023000000;
slave_timing[1][160+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][160+4].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+4].t_rxd1[0][1] = 1728ns;
slave_timing[1][160+4].t_rxd1[1][0] = 1731ns;
slave_timing[1][160+4].t_rxd1[0][2] = 1292ns;
slave_timing[1][160+4].t_rxd1[2][0] = 2087ns;
slave_timing[1][160+4].t_rxd2[0][2] = 1997ns;
slave_timing[1][160+4].t_rxd2[2][0] = 1263ns;
slave_timing[1][160+4].t_rxd2[1][2] = 1650ns;
slave_timing[1][160+4].t_rxd2[2][1] = 1662ns;

slave_timing[1][160+5].info_corner          = 2;
slave_timing[1][160+5].info_temp__j__       = -40;
slave_timing[1][160+5].info_i__quite_rec__  = 0.006000000;
slave_timing[1][160+5].info_dtr__ib__       = -1;
slave_timing[1][160+5].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+5].info_i__max_slave__  = 0.025000000;
slave_timing[1][160+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][160+5].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+5].t_rxd1[0][1] = 1661ns;
slave_timing[1][160+5].t_rxd1[1][0] = 1778ns;
slave_timing[1][160+5].t_rxd1[0][2] = 1270ns;
slave_timing[1][160+5].t_rxd1[2][0] = 2122ns;
slave_timing[1][160+5].t_rxd2[0][2] = 1898ns;
slave_timing[1][160+5].t_rxd2[2][0] = 1346ns;
slave_timing[1][160+5].t_rxd2[1][2] = 1475ns;
slave_timing[1][160+5].t_rxd2[2][1] = 1829ns;

slave_timing[1][160+6].info_corner          = 2;
slave_timing[1][160+6].info_temp__j__       = -40;
slave_timing[1][160+6].info_i__quite_rec__  = 0.006000000;
slave_timing[1][160+6].info_dtr__ib__       = 1;
slave_timing[1][160+6].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+6].info_i__max_slave__  = 0.023000000;
slave_timing[1][160+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][160+6].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+6].t_rxd1[0][1] = 1774ns;
slave_timing[1][160+6].t_rxd1[1][0] = 1687ns;
slave_timing[1][160+6].t_rxd1[0][2] = 1326ns;
slave_timing[1][160+6].t_rxd1[2][0] = 2055ns;
slave_timing[1][160+6].t_rxd2[0][2] = 2121ns;
slave_timing[1][160+6].t_rxd2[2][0] = 1187ns;
slave_timing[1][160+6].t_rxd2[1][2] = 1795ns;
slave_timing[1][160+6].t_rxd2[2][1] = 1534ns;

slave_timing[1][160+7].info_corner          = 2;
slave_timing[1][160+7].info_temp__j__       = -40;
slave_timing[1][160+7].info_i__quite_rec__  = 0.006000000;
slave_timing[1][160+7].info_dtr__ib__       = 1;
slave_timing[1][160+7].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+7].info_i__max_slave__  = 0.025000000;
slave_timing[1][160+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][160+7].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+7].t_rxd1[0][1] = 1701ns;
slave_timing[1][160+7].t_rxd1[1][0] = 1737ns;
slave_timing[1][160+7].t_rxd1[0][2] = 1289ns;
slave_timing[1][160+7].t_rxd1[2][0] = 2090ns;
slave_timing[1][160+7].t_rxd2[0][2] = 1977ns;
slave_timing[1][160+7].t_rxd2[2][0] = 1280ns;
slave_timing[1][160+7].t_rxd2[1][2] = 1600ns;
slave_timing[1][160+7].t_rxd2[2][1] = 1704ns;

slave_timing[1][160+8].info_corner          = 2;
slave_timing[1][160+8].info_temp__j__       = -40;
slave_timing[1][160+8].info_i__quite_rec__  = 0.003000000;
slave_timing[1][160+8].info_dtr__ib__       = -1;
slave_timing[1][160+8].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+8].info_i__max_slave__  = 0.023000000;
slave_timing[1][160+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][160+8].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+8].t_rxd1[0][1] = 1644ns;
slave_timing[1][160+8].t_rxd1[1][0] = 1672ns;
slave_timing[1][160+8].t_rxd1[0][2] = 1239ns;
slave_timing[1][160+8].t_rxd1[2][0] = 2026ns;
slave_timing[1][160+8].t_rxd2[0][2] = 1992ns;
slave_timing[1][160+8].t_rxd2[2][0] = 1251ns;
slave_timing[1][160+8].t_rxd2[1][2] = 1631ns;
slave_timing[1][160+8].t_rxd2[2][1] = 1664ns;

slave_timing[1][160+9].info_corner          = 2;
slave_timing[1][160+9].info_temp__j__       = -40;
slave_timing[1][160+9].info_i__quite_rec__  = 0.003000000;
slave_timing[1][160+9].info_dtr__ib__       = -1;
slave_timing[1][160+9].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+9].info_i__max_slave__  = 0.025000000;
slave_timing[1][160+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][160+9].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+9].t_rxd1[0][1] = 1585ns;
slave_timing[1][160+9].t_rxd1[1][0] = 1719ns;
slave_timing[1][160+9].t_rxd1[0][2] = 1205ns;
slave_timing[1][160+9].t_rxd1[2][0] = 2062ns;
slave_timing[1][160+9].t_rxd2[0][2] = 1873ns;
slave_timing[1][160+9].t_rxd2[2][0] = 1334ns;
slave_timing[1][160+9].t_rxd2[1][2] = 1454ns;
slave_timing[1][160+9].t_rxd2[2][1] = 1835ns;

slave_timing[1][160+10].info_corner          = 2;
slave_timing[1][160+10].info_temp__j__       = -40;
slave_timing[1][160+10].info_i__quite_rec__  = 0.003000000;
slave_timing[1][160+10].info_dtr__ib__       = 1;
slave_timing[1][160+10].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+10].info_i__max_slave__  = 0.023000000;
slave_timing[1][160+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][160+10].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+10].t_rxd1[0][1] = 1697ns;
slave_timing[1][160+10].t_rxd1[1][0] = 1632ns;
slave_timing[1][160+10].t_rxd1[0][2] = 1251ns;
slave_timing[1][160+10].t_rxd1[2][0] = 2000ns;
slave_timing[1][160+10].t_rxd2[0][2] = 2078ns;
slave_timing[1][160+10].t_rxd2[2][0] = 1183ns;
slave_timing[1][160+10].t_rxd2[1][2] = 1777ns;
slave_timing[1][160+10].t_rxd2[2][1] = 1537ns;

slave_timing[1][160+11].info_corner          = 2;
slave_timing[1][160+11].info_temp__j__       = -40;
slave_timing[1][160+11].info_i__quite_rec__  = 0.003000000;
slave_timing[1][160+11].info_dtr__ib__       = 1;
slave_timing[1][160+11].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+11].info_i__max_slave__  = 0.025000000;
slave_timing[1][160+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][160+11].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+11].t_rxd1[0][1] = 1627ns;
slave_timing[1][160+11].t_rxd1[1][0] = 1683ns;
slave_timing[1][160+11].t_rxd1[0][2] = 1228ns;
slave_timing[1][160+11].t_rxd1[2][0] = 2034ns;
slave_timing[1][160+11].t_rxd2[0][2] = 1958ns;
slave_timing[1][160+11].t_rxd2[2][0] = 1273ns;
slave_timing[1][160+11].t_rxd2[1][2] = 1581ns;
slave_timing[1][160+11].t_rxd2[2][1] = 1706ns;

slave_timing[1][160+12].info_corner          = 2;
slave_timing[1][160+12].info_temp__j__       = -40;
slave_timing[1][160+12].info_i__quite_rec__  = 0.003000000;
slave_timing[1][160+12].info_dtr__ib__       = -1;
slave_timing[1][160+12].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+12].info_i__max_slave__  = 0.023000000;
slave_timing[1][160+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][160+12].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+12].t_rxd1[0][1] = 1720ns;
slave_timing[1][160+12].t_rxd1[1][0] = 1740ns;
slave_timing[1][160+12].t_rxd1[0][2] = 1302ns;
slave_timing[1][160+12].t_rxd1[2][0] = 2093ns;
slave_timing[1][160+12].t_rxd2[0][2] = 2007ns;
slave_timing[1][160+12].t_rxd2[2][0] = 1270ns;
slave_timing[1][160+12].t_rxd2[1][2] = 1640ns;
slave_timing[1][160+12].t_rxd2[2][1] = 1652ns;

slave_timing[1][160+13].info_corner          = 2;
slave_timing[1][160+13].info_temp__j__       = -40;
slave_timing[1][160+13].info_i__quite_rec__  = 0.003000000;
slave_timing[1][160+13].info_dtr__ib__       = -1;
slave_timing[1][160+13].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+13].info_i__max_slave__  = 0.025000000;
slave_timing[1][160+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][160+13].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+13].t_rxd1[0][1] = 1656ns;
slave_timing[1][160+13].t_rxd1[1][0] = 1788ns;
slave_timing[1][160+13].t_rxd1[0][2] = 1266ns;
slave_timing[1][160+13].t_rxd1[2][0] = 2126ns;
slave_timing[1][160+13].t_rxd2[0][2] = 1891ns;
slave_timing[1][160+13].t_rxd2[2][0] = 1351ns;
slave_timing[1][160+13].t_rxd2[1][2] = 1468ns;
slave_timing[1][160+13].t_rxd2[2][1] = 1846ns;

slave_timing[1][160+14].info_corner          = 2;
slave_timing[1][160+14].info_temp__j__       = -40;
slave_timing[1][160+14].info_i__quite_rec__  = 0.003000000;
slave_timing[1][160+14].info_dtr__ib__       = 1;
slave_timing[1][160+14].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+14].info_i__max_slave__  = 0.023000000;
slave_timing[1][160+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][160+14].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+14].t_rxd1[0][1] = 1764ns;
slave_timing[1][160+14].t_rxd1[1][0] = 1696ns;
slave_timing[1][160+14].t_rxd1[0][2] = 1322ns;
slave_timing[1][160+14].t_rxd1[2][0] = 2059ns;
slave_timing[1][160+14].t_rxd2[0][2] = 2113ns;
slave_timing[1][160+14].t_rxd2[2][0] = 1196ns;
slave_timing[1][160+14].t_rxd2[1][2] = 1786ns;
slave_timing[1][160+14].t_rxd2[2][1] = 1547ns;

slave_timing[1][160+15].info_corner          = 2;
slave_timing[1][160+15].info_temp__j__       = -40;
slave_timing[1][160+15].info_i__quite_rec__  = 0.003000000;
slave_timing[1][160+15].info_dtr__ib__       = 1;
slave_timing[1][160+15].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+15].info_i__max_slave__  = 0.025000000;
slave_timing[1][160+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][160+15].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+15].t_rxd1[0][1] = 1693ns;
slave_timing[1][160+15].t_rxd1[1][0] = 1747ns;
slave_timing[1][160+15].t_rxd1[0][2] = 1272ns;
slave_timing[1][160+15].t_rxd1[2][0] = 2094ns;
slave_timing[1][160+15].t_rxd2[0][2] = 1958ns;
slave_timing[1][160+15].t_rxd2[2][0] = 1287ns;
slave_timing[1][160+15].t_rxd2[1][2] = 1588ns;
slave_timing[1][160+15].t_rxd2[2][1] = 1714ns;

slave_timing[1][160+16].info_corner          = 2;
slave_timing[1][160+16].info_temp__j__       = -40;
slave_timing[1][160+16].info_i__quite_rec__  = 0.000000000;
slave_timing[1][160+16].info_dtr__ib__       = -1;
slave_timing[1][160+16].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+16].info_i__max_slave__  = 0.023000000;
slave_timing[1][160+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][160+16].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+16].t_rxd1[0][1] = 1662ns;
slave_timing[1][160+16].t_rxd1[1][0] = 1660ns;
slave_timing[1][160+16].t_rxd1[0][2] = 1249ns;
slave_timing[1][160+16].t_rxd1[2][0] = 2020ns;
slave_timing[1][160+16].t_rxd2[0][2] = 2001ns;
slave_timing[1][160+16].t_rxd2[2][0] = 1245ns;
slave_timing[1][160+16].t_rxd2[1][2] = 1642ns;
slave_timing[1][160+16].t_rxd2[2][1] = 1651ns;

slave_timing[1][160+17].info_corner          = 2;
slave_timing[1][160+17].info_temp__j__       = -40;
slave_timing[1][160+17].info_i__quite_rec__  = 0.000000000;
slave_timing[1][160+17].info_dtr__ib__       = -1;
slave_timing[1][160+17].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+17].info_i__max_slave__  = 0.025000000;
slave_timing[1][160+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][160+17].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+17].t_rxd1[0][1] = 1598ns;
slave_timing[1][160+17].t_rxd1[1][0] = 1709ns;
slave_timing[1][160+17].t_rxd1[0][2] = 1215ns;
slave_timing[1][160+17].t_rxd1[2][0] = 2054ns;
slave_timing[1][160+17].t_rxd2[0][2] = 1882ns;
slave_timing[1][160+17].t_rxd2[2][0] = 1328ns;
slave_timing[1][160+17].t_rxd2[1][2] = 1465ns;
slave_timing[1][160+17].t_rxd2[2][1] = 1821ns;

slave_timing[1][160+18].info_corner          = 2;
slave_timing[1][160+18].info_temp__j__       = -40;
slave_timing[1][160+18].info_i__quite_rec__  = 0.000000000;
slave_timing[1][160+18].info_dtr__ib__       = 1;
slave_timing[1][160+18].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+18].info_i__max_slave__  = 0.023000000;
slave_timing[1][160+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][160+18].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+18].t_rxd1[0][1] = 1712ns;
slave_timing[1][160+18].t_rxd1[1][0] = 1619ns;
slave_timing[1][160+18].t_rxd1[0][2] = 1274ns;
slave_timing[1][160+18].t_rxd1[2][0] = 1990ns;
slave_timing[1][160+18].t_rxd2[0][2] = 2112ns;
slave_timing[1][160+18].t_rxd2[2][0] = 1169ns;
slave_timing[1][160+18].t_rxd2[1][2] = 1795ns;
slave_timing[1][160+18].t_rxd2[2][1] = 1516ns;

slave_timing[1][160+19].info_corner          = 2;
slave_timing[1][160+19].info_temp__j__       = -40;
slave_timing[1][160+19].info_i__quite_rec__  = 0.000000000;
slave_timing[1][160+19].info_dtr__ib__       = 1;
slave_timing[1][160+19].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+19].info_i__max_slave__  = 0.025000000;
slave_timing[1][160+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][160+19].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+19].t_rxd1[0][1] = 1643ns;
slave_timing[1][160+19].t_rxd1[1][0] = 1670ns;
slave_timing[1][160+19].t_rxd1[0][2] = 1237ns;
slave_timing[1][160+19].t_rxd1[2][0] = 2026ns;
slave_timing[1][160+19].t_rxd2[0][2] = 1964ns;
slave_timing[1][160+19].t_rxd2[2][0] = 1265ns;
slave_timing[1][160+19].t_rxd2[1][2] = 1596ns;
slave_timing[1][160+19].t_rxd2[2][1] = 1686ns;

slave_timing[1][160+20].info_corner          = 2;
slave_timing[1][160+20].info_temp__j__       = -40;
slave_timing[1][160+20].info_i__quite_rec__  = 0.000000000;
slave_timing[1][160+20].info_dtr__ib__       = -1;
slave_timing[1][160+20].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+20].info_i__max_slave__  = 0.023000000;
slave_timing[1][160+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][160+20].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+20].t_rxd1[0][1] = 1737ns;
slave_timing[1][160+20].t_rxd1[1][0] = 1727ns;
slave_timing[1][160+20].t_rxd1[0][2] = 1310ns;
slave_timing[1][160+20].t_rxd1[2][0] = 2083ns;
slave_timing[1][160+20].t_rxd2[0][2] = 2016ns;
slave_timing[1][160+20].t_rxd2[2][0] = 1259ns;
slave_timing[1][160+20].t_rxd2[1][2] = 1653ns;
slave_timing[1][160+20].t_rxd2[2][1] = 1660ns;

slave_timing[1][160+21].info_corner          = 2;
slave_timing[1][160+21].info_temp__j__       = -40;
slave_timing[1][160+21].info_i__quite_rec__  = 0.000000000;
slave_timing[1][160+21].info_dtr__ib__       = -1;
slave_timing[1][160+21].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+21].info_i__max_slave__  = 0.025000000;
slave_timing[1][160+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][160+21].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+21].t_rxd1[0][1] = 1670ns;
slave_timing[1][160+21].t_rxd1[1][0] = 1775ns;
slave_timing[1][160+21].t_rxd1[0][2] = 1274ns;
slave_timing[1][160+21].t_rxd1[2][0] = 2120ns;
slave_timing[1][160+21].t_rxd2[0][2] = 1897ns;
slave_timing[1][160+21].t_rxd2[2][0] = 1344ns;
slave_timing[1][160+21].t_rxd2[1][2] = 1479ns;
slave_timing[1][160+21].t_rxd2[2][1] = 1831ns;

slave_timing[1][160+22].info_corner          = 2;
slave_timing[1][160+22].info_temp__j__       = -40;
slave_timing[1][160+22].info_i__quite_rec__  = 0.000000000;
slave_timing[1][160+22].info_dtr__ib__       = 1;
slave_timing[1][160+22].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+22].info_i__max_slave__  = 0.023000000;
slave_timing[1][160+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][160+22].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+22].t_rxd1[0][1] = 1780ns;
slave_timing[1][160+22].t_rxd1[1][0] = 1679ns;
slave_timing[1][160+22].t_rxd1[0][2] = 1332ns;
slave_timing[1][160+22].t_rxd1[2][0] = 2052ns;
slave_timing[1][160+22].t_rxd2[0][2] = 2126ns;
slave_timing[1][160+22].t_rxd2[2][0] = 1185ns;
slave_timing[1][160+22].t_rxd2[1][2] = 1804ns;
slave_timing[1][160+22].t_rxd2[2][1] = 1527ns;

slave_timing[1][160+23].info_corner          = 2;
slave_timing[1][160+23].info_temp__j__       = -40;
slave_timing[1][160+23].info_i__quite_rec__  = 0.000000000;
slave_timing[1][160+23].info_dtr__ib__       = 1;
slave_timing[1][160+23].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+23].info_i__max_slave__  = 0.025000000;
slave_timing[1][160+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][160+23].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+23].t_rxd1[0][1] = 1709ns;
slave_timing[1][160+23].t_rxd1[1][0] = 1733ns;
slave_timing[1][160+23].t_rxd1[0][2] = 1294ns;
slave_timing[1][160+23].t_rxd1[2][0] = 2087ns;
slave_timing[1][160+23].t_rxd2[0][2] = 1979ns;
slave_timing[1][160+23].t_rxd2[2][0] = 1275ns;
slave_timing[1][160+23].t_rxd2[1][2] = 1606ns;
slave_timing[1][160+23].t_rxd2[2][1] = 1695ns;

slave_timing[1][160+24].info_corner          = 2;
slave_timing[1][160+24].info_temp__j__       = -40;
slave_timing[1][160+24].info_i__quite_rec__  = 0.040000000;
slave_timing[1][160+24].info_dtr__ib__       = -1;
slave_timing[1][160+24].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+24].info_i__max_slave__  = 0.023000000;
slave_timing[1][160+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][160+24].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+24].t_rxd1[0][1] = 1656ns;
slave_timing[1][160+24].t_rxd1[1][0] = 1650ns;
slave_timing[1][160+24].t_rxd1[0][2] = 1244ns;
slave_timing[1][160+24].t_rxd1[2][0] = 2011ns;
slave_timing[1][160+24].t_rxd2[0][2] = 2001ns;
slave_timing[1][160+24].t_rxd2[2][0] = 1243ns;
slave_timing[1][160+24].t_rxd2[1][2] = 1644ns;
slave_timing[1][160+24].t_rxd2[2][1] = 1647ns;

slave_timing[1][160+25].info_corner          = 2;
slave_timing[1][160+25].info_temp__j__       = -40;
slave_timing[1][160+25].info_i__quite_rec__  = 0.040000000;
slave_timing[1][160+25].info_dtr__ib__       = -1;
slave_timing[1][160+25].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+25].info_i__max_slave__  = 0.025000000;
slave_timing[1][160+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][160+25].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+25].t_rxd1[0][1] = 1589ns;
slave_timing[1][160+25].t_rxd1[1][0] = 1701ns;
slave_timing[1][160+25].t_rxd1[0][2] = 1208ns;
slave_timing[1][160+25].t_rxd1[2][0] = 2046ns;
slave_timing[1][160+25].t_rxd2[0][2] = 1881ns;
slave_timing[1][160+25].t_rxd2[2][0] = 1327ns;
slave_timing[1][160+25].t_rxd2[1][2] = 1470ns;
slave_timing[1][160+25].t_rxd2[2][1] = 1819ns;

slave_timing[1][160+26].info_corner          = 2;
slave_timing[1][160+26].info_temp__j__       = -40;
slave_timing[1][160+26].info_i__quite_rec__  = 0.040000000;
slave_timing[1][160+26].info_dtr__ib__       = 1;
slave_timing[1][160+26].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+26].info_i__max_slave__  = 0.023000000;
slave_timing[1][160+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][160+26].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+26].t_rxd1[0][1] = 1696ns;
slave_timing[1][160+26].t_rxd1[1][0] = 1624ns;
slave_timing[1][160+26].t_rxd1[0][2] = 1263ns;
slave_timing[1][160+26].t_rxd1[2][0] = 1992ns;
slave_timing[1][160+26].t_rxd2[0][2] = 2105ns;
slave_timing[1][160+26].t_rxd2[2][0] = 1175ns;
slave_timing[1][160+26].t_rxd2[1][2] = 1783ns;
slave_timing[1][160+26].t_rxd2[2][1] = 1525ns;

slave_timing[1][160+27].info_corner          = 2;
slave_timing[1][160+27].info_temp__j__       = -40;
slave_timing[1][160+27].info_i__quite_rec__  = 0.040000000;
slave_timing[1][160+27].info_dtr__ib__       = 1;
slave_timing[1][160+27].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+27].info_i__max_slave__  = 0.025000000;
slave_timing[1][160+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][160+27].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+27].t_rxd1[0][1] = 1625ns;
slave_timing[1][160+27].t_rxd1[1][0] = 1673ns;
slave_timing[1][160+27].t_rxd1[0][2] = 1216ns;
slave_timing[1][160+27].t_rxd1[2][0] = 2026ns;
slave_timing[1][160+27].t_rxd2[0][2] = 1944ns;
slave_timing[1][160+27].t_rxd2[2][0] = 1266ns;
slave_timing[1][160+27].t_rxd2[1][2] = 1586ns;
slave_timing[1][160+27].t_rxd2[2][1] = 1697ns;

slave_timing[1][160+28].info_corner          = 2;
slave_timing[1][160+28].info_temp__j__       = -40;
slave_timing[1][160+28].info_i__quite_rec__  = 0.040000000;
slave_timing[1][160+28].info_dtr__ib__       = -1;
slave_timing[1][160+28].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+28].info_i__max_slave__  = 0.023000000;
slave_timing[1][160+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][160+28].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+28].t_rxd1[0][1] = 1695ns;
slave_timing[1][160+28].t_rxd1[1][0] = 1689ns;
slave_timing[1][160+28].t_rxd1[0][2] = 1281ns;
slave_timing[1][160+28].t_rxd1[2][0] = 2047ns;
slave_timing[1][160+28].t_rxd2[0][2] = 2012ns;
slave_timing[1][160+28].t_rxd2[2][0] = 1259ns;
slave_timing[1][160+28].t_rxd2[1][2] = 1656ns;
slave_timing[1][160+28].t_rxd2[2][1] = 1657ns;

slave_timing[1][160+29].info_corner          = 2;
slave_timing[1][160+29].info_temp__j__       = -40;
slave_timing[1][160+29].info_i__quite_rec__  = 0.040000000;
slave_timing[1][160+29].info_dtr__ib__       = -1;
slave_timing[1][160+29].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+29].info_i__max_slave__  = 0.025000000;
slave_timing[1][160+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][160+29].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+29].t_rxd1[0][1] = 1629ns;
slave_timing[1][160+29].t_rxd1[1][0] = 1738ns;
slave_timing[1][160+29].t_rxd1[0][2] = 1244ns;
slave_timing[1][160+29].t_rxd1[2][0] = 2083ns;
slave_timing[1][160+29].t_rxd2[0][2] = 1894ns;
slave_timing[1][160+29].t_rxd2[2][0] = 1341ns;
slave_timing[1][160+29].t_rxd2[1][2] = 1484ns;
slave_timing[1][160+29].t_rxd2[2][1] = 1827ns;

slave_timing[1][160+30].info_corner          = 2;
slave_timing[1][160+30].info_temp__j__       = -40;
slave_timing[1][160+30].info_i__quite_rec__  = 0.040000000;
slave_timing[1][160+30].info_dtr__ib__       = 1;
slave_timing[1][160+30].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+30].info_i__max_slave__  = 0.023000000;
slave_timing[1][160+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][160+30].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+30].t_rxd1[0][1] = 1732ns;
slave_timing[1][160+30].t_rxd1[1][0] = 1661ns;
slave_timing[1][160+30].t_rxd1[0][2] = 1298ns;
slave_timing[1][160+30].t_rxd1[2][0] = 2026ns;
slave_timing[1][160+30].t_rxd2[0][2] = 2113ns;
slave_timing[1][160+30].t_rxd2[2][0] = 1190ns;
slave_timing[1][160+30].t_rxd2[1][2] = 1795ns;
slave_timing[1][160+30].t_rxd2[2][1] = 1537ns;

slave_timing[1][160+31].info_corner          = 2;
slave_timing[1][160+31].info_temp__j__       = -40;
slave_timing[1][160+31].info_i__quite_rec__  = 0.040000000;
slave_timing[1][160+31].info_dtr__ib__       = 1;
slave_timing[1][160+31].info_i__offset_rec__ = 0.000000000;
slave_timing[1][160+31].info_i__max_slave__  = 0.025000000;
slave_timing[1][160+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][160+31].info_r__dsi_bus__    = 5.000;

slave_timing[1][160+31].t_rxd1[0][1] = 1664ns;
slave_timing[1][160+31].t_rxd1[1][0] = 1706ns;
slave_timing[1][160+31].t_rxd1[0][2] = 1260ns;
slave_timing[1][160+31].t_rxd1[2][0] = 2060ns;
slave_timing[1][160+31].t_rxd2[0][2] = 1971ns;
slave_timing[1][160+31].t_rxd2[2][0] = 1282ns;
slave_timing[1][160+31].t_rxd2[1][2] = 1600ns;
slave_timing[1][160+31].t_rxd2[2][1] = 1702ns;

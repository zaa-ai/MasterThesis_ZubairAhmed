/* ###   interface instances   ###################################################### */

OTP_test_registers_OTP_WRITE_PULSE_WIDTH_if OTP_test_registers_OTP_WRITE_PULSE_WIDTH (); 


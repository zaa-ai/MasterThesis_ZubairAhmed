
slave_timing[3][0].info_corner          = 0;
slave_timing[3][0].info_temp__j__       = 25;
slave_timing[3][0].info_i__quite_rec__  = 0.006000000;
slave_timing[3][0].info_dtr__ib__       = -1;
slave_timing[3][0].info_i__offset_rec__ = -0.001000000;
slave_timing[3][0].info_i__max_slave__  = 0.021000000;
slave_timing[3][0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][0].info_r__dsi_bus__    = 5.000;

slave_timing[3][0].t_rxd1[0][1] = 3536ns;
slave_timing[3][0].t_rxd1[1][0] = 2520ns;
slave_timing[3][0].t_rxd1[0][2] = 2426ns;
slave_timing[3][0].t_rxd1[2][0] = 3218ns;
slave_timing[3][0].t_rxd2[0][2] = 3940ns;
slave_timing[3][0].t_rxd2[2][0] = 1943ns;
slave_timing[3][0].t_rxd2[1][2] = 3565ns;
slave_timing[3][0].t_rxd2[2][1] = 2525ns;

slave_timing[3][1].info_corner          = 0;
slave_timing[3][1].info_temp__j__       = 25;
slave_timing[3][1].info_i__quite_rec__  = 0.006000000;
slave_timing[3][1].info_dtr__ib__       = -1;
slave_timing[3][1].info_i__offset_rec__ = 0.001000000;
slave_timing[3][1].info_i__max_slave__  = 0.021000000;
slave_timing[3][1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][1].info_r__dsi_bus__    = 5.000;

slave_timing[3][1].t_rxd1[0][1] = 2964ns;
slave_timing[3][1].t_rxd1[1][0] = 2976ns;
slave_timing[3][1].t_rxd1[0][2] = 2190ns;
slave_timing[3][1].t_rxd1[2][0] = 3515ns;
slave_timing[3][1].t_rxd2[0][2] = 3520ns;
slave_timing[3][1].t_rxd2[2][0] = 2208ns;
slave_timing[3][1].t_rxd2[1][2] = 2987ns;
slave_timing[3][1].t_rxd2[2][1] = 2982ns;

slave_timing[3][2].info_corner          = 0;
slave_timing[3][2].info_temp__j__       = 25;
slave_timing[3][2].info_i__quite_rec__  = 0.006000000;
slave_timing[3][2].info_dtr__ib__       = -1;
slave_timing[3][2].info_i__offset_rec__ = -0.001000000;
slave_timing[3][2].info_i__max_slave__  = 0.027000000;
slave_timing[3][2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][2].info_r__dsi_bus__    = 5.000;

slave_timing[3][2].t_rxd1[0][1] = 2988ns;
slave_timing[3][2].t_rxd1[1][0] = 2797ns;
slave_timing[3][2].t_rxd1[0][2] = 2200ns;
slave_timing[3][2].t_rxd1[2][0] = 3398ns;
slave_timing[3][2].t_rxd2[0][2] = 3175ns;
slave_timing[3][2].t_rxd2[2][0] = 2394ns;
slave_timing[3][2].t_rxd2[1][2] = 2474ns;
slave_timing[3][2].t_rxd2[2][1] = 3419ns;

slave_timing[3][3].info_corner          = 0;
slave_timing[3][3].info_temp__j__       = 25;
slave_timing[3][3].info_i__quite_rec__  = 0.006000000;
slave_timing[3][3].info_dtr__ib__       = -1;
slave_timing[3][3].info_i__offset_rec__ = 0.001000000;
slave_timing[3][3].info_i__max_slave__  = 0.027000000;
slave_timing[3][3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][3].info_r__dsi_bus__    = 5.000;

slave_timing[3][3].t_rxd1[0][1] = 2663ns;
slave_timing[3][3].t_rxd1[1][0] = 3142ns;
slave_timing[3][3].t_rxd1[0][2] = 2016ns;
slave_timing[3][3].t_rxd1[2][0] = 3634ns;
slave_timing[3][3].t_rxd2[0][2] = 2991ns;
slave_timing[3][3].t_rxd2[2][0] = 2547ns;
slave_timing[3][3].t_rxd2[1][2] = 2143ns;
slave_timing[3][3].t_rxd2[2][1] = 3978ns;

slave_timing[3][4].info_corner          = 0;
slave_timing[3][4].info_temp__j__       = 25;
slave_timing[3][4].info_i__quite_rec__  = 0.006000000;
slave_timing[3][4].info_dtr__ib__       = 1;
slave_timing[3][4].info_i__offset_rec__ = -0.001000000;
slave_timing[3][4].info_i__max_slave__  = 0.021000000;
slave_timing[3][4].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][4].info_r__dsi_bus__    = 5.000;

slave_timing[3][4].t_rxd1[0][1] = 3706ns;
slave_timing[3][4].t_rxd1[1][0] = 2453ns;
slave_timing[3][4].t_rxd1[0][2] = 2476ns;
slave_timing[3][4].t_rxd1[2][0] = 3175ns;
slave_timing[3][4].t_rxd2[0][2] = 4353ns;
slave_timing[3][4].t_rxd2[2][0] = 1789ns;
slave_timing[3][4].t_rxd2[1][2] = 4103ns;
slave_timing[3][4].t_rxd2[2][1] = 2302ns;

slave_timing[3][5].info_corner          = 0;
slave_timing[3][5].info_temp__j__       = 25;
slave_timing[3][5].info_i__quite_rec__  = 0.006000000;
slave_timing[3][5].info_dtr__ib__       = 1;
slave_timing[3][5].info_i__offset_rec__ = 0.001000000;
slave_timing[3][5].info_i__max_slave__  = 0.021000000;
slave_timing[3][5].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][5].info_r__dsi_bus__    = 5.000;

slave_timing[3][5].t_rxd1[0][1] = 3080ns;
slave_timing[3][5].t_rxd1[1][0] = 2906ns;
slave_timing[3][5].t_rxd1[0][2] = 2250ns;
slave_timing[3][5].t_rxd1[2][0] = 3469ns;
slave_timing[3][5].t_rxd2[0][2] = 3737ns;
slave_timing[3][5].t_rxd2[2][0] = 2083ns;
slave_timing[3][5].t_rxd2[1][2] = 3296ns;
slave_timing[3][5].t_rxd2[2][1] = 2751ns;

slave_timing[3][6].info_corner          = 0;
slave_timing[3][6].info_temp__j__       = 25;
slave_timing[3][6].info_i__quite_rec__  = 0.006000000;
slave_timing[3][6].info_dtr__ib__       = 1;
slave_timing[3][6].info_i__offset_rec__ = -0.001000000;
slave_timing[3][6].info_i__max_slave__  = 0.027000000;
slave_timing[3][6].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][6].info_r__dsi_bus__    = 5.000;

slave_timing[3][6].t_rxd1[0][1] = 3079ns;
slave_timing[3][6].t_rxd1[1][0] = 2749ns;
slave_timing[3][6].t_rxd1[0][2] = 2244ns;
slave_timing[3][6].t_rxd1[2][0] = 3360ns;
slave_timing[3][6].t_rxd2[0][2] = 3300ns;
slave_timing[3][6].t_rxd2[2][0] = 2302ns;
slave_timing[3][6].t_rxd2[1][2] = 2668ns;
slave_timing[3][6].t_rxd2[2][1] = 3193ns;

slave_timing[3][7].info_corner          = 0;
slave_timing[3][7].info_temp__j__       = 25;
slave_timing[3][7].info_i__quite_rec__  = 0.006000000;
slave_timing[3][7].info_dtr__ib__       = 1;
slave_timing[3][7].info_i__offset_rec__ = 0.001000000;
slave_timing[3][7].info_i__max_slave__  = 0.027000000;
slave_timing[3][7].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][7].info_r__dsi_bus__    = 5.000;

slave_timing[3][7].t_rxd1[0][1] = 2747ns;
slave_timing[3][7].t_rxd1[1][0] = 3082ns;
slave_timing[3][7].t_rxd1[0][2] = 2046ns;
slave_timing[3][7].t_rxd1[2][0] = 3590ns;
slave_timing[3][7].t_rxd2[0][2] = 3087ns;
slave_timing[3][7].t_rxd2[2][0] = 2461ns;
slave_timing[3][7].t_rxd2[1][2] = 2358ns;
slave_timing[3][7].t_rxd2[2][1] = 3633ns;

slave_timing[3][8].info_corner          = 0;
slave_timing[3][8].info_temp__j__       = 25;
slave_timing[3][8].info_i__quite_rec__  = 0.006000000;
slave_timing[3][8].info_dtr__ib__       = -1;
slave_timing[3][8].info_i__offset_rec__ = -0.001000000;
slave_timing[3][8].info_i__max_slave__  = 0.021000000;
slave_timing[3][8].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][8].info_r__dsi_bus__    = 5.000;

slave_timing[3][8].t_rxd1[0][1] = 3774ns;
slave_timing[3][8].t_rxd1[1][0] = 2728ns;
slave_timing[3][8].t_rxd1[0][2] = 2628ns;
slave_timing[3][8].t_rxd1[2][0] = 3448ns;
slave_timing[3][8].t_rxd2[0][2] = 4205ns;
slave_timing[3][8].t_rxd2[2][0] = 2132ns;
slave_timing[3][8].t_rxd2[1][2] = 3807ns;
slave_timing[3][8].t_rxd2[2][1] = 2734ns;

slave_timing[3][9].info_corner          = 0;
slave_timing[3][9].info_temp__j__       = 25;
slave_timing[3][9].info_i__quite_rec__  = 0.006000000;
slave_timing[3][9].info_dtr__ib__       = -1;
slave_timing[3][9].info_i__offset_rec__ = 0.001000000;
slave_timing[3][9].info_i__max_slave__  = 0.021000000;
slave_timing[3][9].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][9].info_r__dsi_bus__    = 5.000;

slave_timing[3][9].t_rxd1[0][1] = 3188ns;
slave_timing[3][9].t_rxd1[1][0] = 3198ns;
slave_timing[3][9].t_rxd1[0][2] = 2384ns;
slave_timing[3][9].t_rxd1[2][0] = 3762ns;
slave_timing[3][9].t_rxd2[0][2] = 3762ns;
slave_timing[3][9].t_rxd2[2][0] = 2402ns;
slave_timing[3][9].t_rxd2[1][2] = 3213ns;
slave_timing[3][9].t_rxd2[2][1] = 3209ns;

slave_timing[3][10].info_corner          = 0;
slave_timing[3][10].info_temp__j__       = 25;
slave_timing[3][10].info_i__quite_rec__  = 0.006000000;
slave_timing[3][10].info_dtr__ib__       = -1;
slave_timing[3][10].info_i__offset_rec__ = -0.001000000;
slave_timing[3][10].info_i__max_slave__  = 0.027000000;
slave_timing[3][10].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][10].info_r__dsi_bus__    = 5.000;

slave_timing[3][10].t_rxd1[0][1] = 3215ns;
slave_timing[3][10].t_rxd1[1][0] = 3018ns;
slave_timing[3][10].t_rxd1[0][2] = 2395ns;
slave_timing[3][10].t_rxd1[2][0] = 3634ns;
slave_timing[3][10].t_rxd2[0][2] = 3404ns;
slave_timing[3][10].t_rxd2[2][0] = 2589ns;
slave_timing[3][10].t_rxd2[1][2] = 2673ns;
slave_timing[3][10].t_rxd2[2][1] = 3658ns;

slave_timing[3][11].info_corner          = 0;
slave_timing[3][11].info_temp__j__       = 25;
slave_timing[3][11].info_i__quite_rec__  = 0.006000000;
slave_timing[3][11].info_dtr__ib__       = -1;
slave_timing[3][11].info_i__offset_rec__ = 0.001000000;
slave_timing[3][11].info_i__max_slave__  = 0.027000000;
slave_timing[3][11].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][11].info_r__dsi_bus__    = 5.000;

slave_timing[3][11].t_rxd1[0][1] = 2839ns;
slave_timing[3][11].t_rxd1[1][0] = 3415ns;
slave_timing[3][11].t_rxd1[0][2] = 2187ns;
slave_timing[3][11].t_rxd1[2][0] = 3913ns;
slave_timing[3][11].t_rxd2[0][2] = 3197ns;
slave_timing[3][11].t_rxd2[2][0] = 2774ns;
slave_timing[3][11].t_rxd2[1][2] = 2297ns;
slave_timing[3][11].t_rxd2[2][1] = 4370ns;

slave_timing[3][12].info_corner          = 0;
slave_timing[3][12].info_temp__j__       = 25;
slave_timing[3][12].info_i__quite_rec__  = 0.006000000;
slave_timing[3][12].info_dtr__ib__       = 1;
slave_timing[3][12].info_i__offset_rec__ = -0.001000000;
slave_timing[3][12].info_i__max_slave__  = 0.021000000;
slave_timing[3][12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][12].info_r__dsi_bus__    = 5.000;

slave_timing[3][12].t_rxd1[0][1] = 3961ns;
slave_timing[3][12].t_rxd1[1][0] = 2657ns;
slave_timing[3][12].t_rxd1[0][2] = 2684ns;
slave_timing[3][12].t_rxd1[2][0] = 3405ns;
slave_timing[3][12].t_rxd2[0][2] = 4655ns;
slave_timing[3][12].t_rxd2[2][0] = 1977ns;
slave_timing[3][12].t_rxd2[1][2] = 4368ns;
slave_timing[3][12].t_rxd2[2][1] = 2500ns;

slave_timing[3][13].info_corner          = 0;
slave_timing[3][13].info_temp__j__       = 25;
slave_timing[3][13].info_i__quite_rec__  = 0.006000000;
slave_timing[3][13].info_dtr__ib__       = 1;
slave_timing[3][13].info_i__offset_rec__ = 0.001000000;
slave_timing[3][13].info_i__max_slave__  = 0.021000000;
slave_timing[3][13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][13].info_r__dsi_bus__    = 5.000;

slave_timing[3][13].t_rxd1[0][1] = 3310ns;
slave_timing[3][13].t_rxd1[1][0] = 3128ns;
slave_timing[3][13].t_rxd1[0][2] = 2441ns;
slave_timing[3][13].t_rxd1[2][0] = 3709ns;
slave_timing[3][13].t_rxd2[0][2] = 3991ns;
slave_timing[3][13].t_rxd2[2][0] = 2274ns;
slave_timing[3][13].t_rxd2[1][2] = 3531ns;
slave_timing[3][13].t_rxd2[2][1] = 2968ns;

slave_timing[3][14].info_corner          = 0;
slave_timing[3][14].info_temp__j__       = 25;
slave_timing[3][14].info_i__quite_rec__  = 0.006000000;
slave_timing[3][14].info_dtr__ib__       = 1;
slave_timing[3][14].info_i__offset_rec__ = -0.001000000;
slave_timing[3][14].info_i__max_slave__  = 0.027000000;
slave_timing[3][14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][14].info_r__dsi_bus__    = 5.000;

slave_timing[3][14].t_rxd1[0][1] = 3304ns;
slave_timing[3][14].t_rxd1[1][0] = 2964ns;
slave_timing[3][14].t_rxd1[0][2] = 2443ns;
slave_timing[3][14].t_rxd1[2][0] = 3598ns;
slave_timing[3][14].t_rxd2[0][2] = 3538ns;
slave_timing[3][14].t_rxd2[2][0] = 2501ns;
slave_timing[3][14].t_rxd2[1][2] = 2885ns;
slave_timing[3][14].t_rxd2[2][1] = 3426ns;

slave_timing[3][15].info_corner          = 0;
slave_timing[3][15].info_temp__j__       = 25;
slave_timing[3][15].info_i__quite_rec__  = 0.006000000;
slave_timing[3][15].info_dtr__ib__       = 1;
slave_timing[3][15].info_i__offset_rec__ = 0.001000000;
slave_timing[3][15].info_i__max_slave__  = 0.027000000;
slave_timing[3][15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][15].info_r__dsi_bus__    = 5.000;

slave_timing[3][15].t_rxd1[0][1] = 2959ns;
slave_timing[3][15].t_rxd1[1][0] = 3311ns;
slave_timing[3][15].t_rxd1[0][2] = 2260ns;
slave_timing[3][15].t_rxd1[2][0] = 3836ns;
slave_timing[3][15].t_rxd2[0][2] = 3337ns;
slave_timing[3][15].t_rxd2[2][0] = 2667ns;
slave_timing[3][15].t_rxd2[1][2] = 2561ns;
slave_timing[3][15].t_rxd2[2][1] = 3881ns;

slave_timing[3][16].info_corner          = 0;
slave_timing[3][16].info_temp__j__       = 25;
slave_timing[3][16].info_i__quite_rec__  = 0.003000000;
slave_timing[3][16].info_dtr__ib__       = -1;
slave_timing[3][16].info_i__offset_rec__ = -0.001000000;
slave_timing[3][16].info_i__max_slave__  = 0.021000000;
slave_timing[3][16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][16].info_r__dsi_bus__    = 5.000;

slave_timing[3][16].t_rxd1[0][1] = 3497ns;
slave_timing[3][16].t_rxd1[1][0] = 2535ns;
slave_timing[3][16].t_rxd1[0][2] = 2417ns;
slave_timing[3][16].t_rxd1[2][0] = 3224ns;
slave_timing[3][16].t_rxd2[0][2] = 3915ns;
slave_timing[3][16].t_rxd2[2][0] = 1954ns;
slave_timing[3][16].t_rxd2[1][2] = 3533ns;
slave_timing[3][16].t_rxd2[2][1] = 2541ns;

slave_timing[3][17].info_corner          = 0;
slave_timing[3][17].info_temp__j__       = 25;
slave_timing[3][17].info_i__quite_rec__  = 0.003000000;
slave_timing[3][17].info_dtr__ib__       = -1;
slave_timing[3][17].info_i__offset_rec__ = 0.001000000;
slave_timing[3][17].info_i__max_slave__  = 0.021000000;
slave_timing[3][17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][17].info_r__dsi_bus__    = 5.000;

slave_timing[3][17].t_rxd1[0][1] = 2990ns;
slave_timing[3][17].t_rxd1[1][0] = 2947ns;
slave_timing[3][17].t_rxd1[0][2] = 2179ns;
slave_timing[3][17].t_rxd1[2][0] = 3495ns;
slave_timing[3][17].t_rxd2[0][2] = 3503ns;
slave_timing[3][17].t_rxd2[2][0] = 2195ns;
slave_timing[3][17].t_rxd2[1][2] = 3014ns;
slave_timing[3][17].t_rxd2[2][1] = 2954ns;

slave_timing[3][18].info_corner          = 0;
slave_timing[3][18].info_temp__j__       = 25;
slave_timing[3][18].info_i__quite_rec__  = 0.003000000;
slave_timing[3][18].info_dtr__ib__       = -1;
slave_timing[3][18].info_i__offset_rec__ = -0.001000000;
slave_timing[3][18].info_i__max_slave__  = 0.027000000;
slave_timing[3][18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][18].info_r__dsi_bus__    = 5.000;

slave_timing[3][18].t_rxd1[0][1] = 3007ns;
slave_timing[3][18].t_rxd1[1][0] = 2777ns;
slave_timing[3][18].t_rxd1[0][2] = 2208ns;
slave_timing[3][18].t_rxd1[2][0] = 3378ns;
slave_timing[3][18].t_rxd2[0][2] = 3181ns;
slave_timing[3][18].t_rxd2[2][0] = 2380ns;
slave_timing[3][18].t_rxd2[1][2] = 2489ns;
slave_timing[3][18].t_rxd2[2][1] = 3389ns;

slave_timing[3][19].info_corner          = 0;
slave_timing[3][19].info_temp__j__       = 25;
slave_timing[3][19].info_i__quite_rec__  = 0.003000000;
slave_timing[3][19].info_dtr__ib__       = -1;
slave_timing[3][19].info_i__offset_rec__ = 0.001000000;
slave_timing[3][19].info_i__max_slave__  = 0.027000000;
slave_timing[3][19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][19].info_r__dsi_bus__    = 5.000;

slave_timing[3][19].t_rxd1[0][1] = 2648ns;
slave_timing[3][19].t_rxd1[1][0] = 3157ns;
slave_timing[3][19].t_rxd1[0][2] = 2009ns;
slave_timing[3][19].t_rxd1[2][0] = 3645ns;
slave_timing[3][19].t_rxd2[0][2] = 2981ns;
slave_timing[3][19].t_rxd2[2][0] = 2553ns;
slave_timing[3][19].t_rxd2[1][2] = 2127ns;
slave_timing[3][19].t_rxd2[2][1] = 4014ns;

slave_timing[3][20].info_corner          = 0;
slave_timing[3][20].info_temp__j__       = 25;
slave_timing[3][20].info_i__quite_rec__  = 0.003000000;
slave_timing[3][20].info_dtr__ib__       = 1;
slave_timing[3][20].info_i__offset_rec__ = -0.001000000;
slave_timing[3][20].info_i__max_slave__  = 0.021000000;
slave_timing[3][20].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][20].info_r__dsi_bus__    = 5.000;

slave_timing[3][20].t_rxd1[0][1] = 3668ns;
slave_timing[3][20].t_rxd1[1][0] = 2471ns;
slave_timing[3][20].t_rxd1[0][2] = 2466ns;
slave_timing[3][20].t_rxd1[2][0] = 3183ns;
slave_timing[3][20].t_rxd2[0][2] = 4321ns;
slave_timing[3][20].t_rxd2[2][0] = 1802ns;
slave_timing[3][20].t_rxd2[1][2] = 4055ns;
slave_timing[3][20].t_rxd2[2][1] = 2314ns;

slave_timing[3][21].info_corner          = 0;
slave_timing[3][21].info_temp__j__       = 25;
slave_timing[3][21].info_i__quite_rec__  = 0.003000000;
slave_timing[3][21].info_dtr__ib__       = 1;
slave_timing[3][21].info_i__offset_rec__ = 0.001000000;
slave_timing[3][21].info_i__max_slave__  = 0.021000000;
slave_timing[3][21].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][21].info_r__dsi_bus__    = 5.000;

slave_timing[3][21].t_rxd1[0][1] = 3061ns;
slave_timing[3][21].t_rxd1[1][0] = 2920ns;
slave_timing[3][21].t_rxd1[0][2] = 2238ns;
slave_timing[3][21].t_rxd1[2][0] = 3477ns;
slave_timing[3][21].t_rxd2[0][2] = 3720ns;
slave_timing[3][21].t_rxd2[2][0] = 2093ns;
slave_timing[3][21].t_rxd2[1][2] = 3269ns;
slave_timing[3][21].t_rxd2[2][1] = 2769ns;

slave_timing[3][22].info_corner          = 0;
slave_timing[3][22].info_temp__j__       = 25;
slave_timing[3][22].info_i__quite_rec__  = 0.003000000;
slave_timing[3][22].info_dtr__ib__       = 1;
slave_timing[3][22].info_i__offset_rec__ = -0.001000000;
slave_timing[3][22].info_i__max_slave__  = 0.027000000;
slave_timing[3][22].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][22].info_r__dsi_bus__    = 5.000;

slave_timing[3][22].t_rxd1[0][1] = 3063ns;
slave_timing[3][22].t_rxd1[1][0] = 2757ns;
slave_timing[3][22].t_rxd1[0][2] = 2238ns;
slave_timing[3][22].t_rxd1[2][0] = 3364ns;
slave_timing[3][22].t_rxd2[0][2] = 3288ns;
slave_timing[3][22].t_rxd2[2][0] = 2309ns;
slave_timing[3][22].t_rxd2[1][2] = 2656ns;
slave_timing[3][22].t_rxd2[2][1] = 3200ns;

slave_timing[3][23].info_corner          = 0;
slave_timing[3][23].info_temp__j__       = 25;
slave_timing[3][23].info_i__quite_rec__  = 0.003000000;
slave_timing[3][23].info_dtr__ib__       = 1;
slave_timing[3][23].info_i__offset_rec__ = 0.001000000;
slave_timing[3][23].info_i__max_slave__  = 0.027000000;
slave_timing[3][23].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][23].info_r__dsi_bus__    = 5.000;

slave_timing[3][23].t_rxd1[0][1] = 2733ns;
slave_timing[3][23].t_rxd1[1][0] = 3091ns;
slave_timing[3][23].t_rxd1[0][2] = 2060ns;
slave_timing[3][23].t_rxd1[2][0] = 3596ns;
slave_timing[3][23].t_rxd2[0][2] = 3095ns;
slave_timing[3][23].t_rxd2[2][0] = 2467ns;
slave_timing[3][23].t_rxd2[1][2] = 2342ns;
slave_timing[3][23].t_rxd2[2][1] = 3650ns;

slave_timing[3][24].info_corner          = 0;
slave_timing[3][24].info_temp__j__       = 25;
slave_timing[3][24].info_i__quite_rec__  = 0.003000000;
slave_timing[3][24].info_dtr__ib__       = -1;
slave_timing[3][24].info_i__offset_rec__ = -0.001000000;
slave_timing[3][24].info_i__max_slave__  = 0.021000000;
slave_timing[3][24].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][24].info_r__dsi_bus__    = 5.000;

slave_timing[3][24].t_rxd1[0][1] = 3743ns;
slave_timing[3][24].t_rxd1[1][0] = 2741ns;
slave_timing[3][24].t_rxd1[0][2] = 2619ns;
slave_timing[3][24].t_rxd1[2][0] = 3456ns;
slave_timing[3][24].t_rxd2[0][2] = 4183ns;
slave_timing[3][24].t_rxd2[2][0] = 2143ns;
slave_timing[3][24].t_rxd2[1][2] = 3776ns;
slave_timing[3][24].t_rxd2[2][1] = 2751ns;

slave_timing[3][25].info_corner          = 0;
slave_timing[3][25].info_temp__j__       = 25;
slave_timing[3][25].info_i__quite_rec__  = 0.003000000;
slave_timing[3][25].info_dtr__ib__       = -1;
slave_timing[3][25].info_i__offset_rec__ = 0.001000000;
slave_timing[3][25].info_i__max_slave__  = 0.021000000;
slave_timing[3][25].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][25].info_r__dsi_bus__    = 5.000;

slave_timing[3][25].t_rxd1[0][1] = 3168ns;
slave_timing[3][25].t_rxd1[1][0] = 3214ns;
slave_timing[3][25].t_rxd1[0][2] = 2375ns;
slave_timing[3][25].t_rxd1[2][0] = 3771ns;
slave_timing[3][25].t_rxd2[0][2] = 3747ns;
slave_timing[3][25].t_rxd2[2][0] = 2413ns;
slave_timing[3][25].t_rxd2[1][2] = 3192ns;
slave_timing[3][25].t_rxd2[2][1] = 3224ns;

slave_timing[3][26].info_corner          = 0;
slave_timing[3][26].info_temp__j__       = 25;
slave_timing[3][26].info_i__quite_rec__  = 0.003000000;
slave_timing[3][26].info_dtr__ib__       = -1;
slave_timing[3][26].info_i__offset_rec__ = -0.001000000;
slave_timing[3][26].info_i__max_slave__  = 0.027000000;
slave_timing[3][26].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][26].info_r__dsi_bus__    = 5.000;

slave_timing[3][26].t_rxd1[0][1] = 3195ns;
slave_timing[3][26].t_rxd1[1][0] = 3027ns;
slave_timing[3][26].t_rxd1[0][2] = 2406ns;
slave_timing[3][26].t_rxd1[2][0] = 3617ns;
slave_timing[3][26].t_rxd2[0][2] = 3417ns;
slave_timing[3][26].t_rxd2[2][0] = 2582ns;
slave_timing[3][26].t_rxd2[1][2] = 2665ns;
slave_timing[3][26].t_rxd2[2][1] = 3674ns;

slave_timing[3][27].info_corner          = 0;
slave_timing[3][27].info_temp__j__       = 25;
slave_timing[3][27].info_i__quite_rec__  = 0.003000000;
slave_timing[3][27].info_dtr__ib__       = -1;
slave_timing[3][27].info_i__offset_rec__ = 0.001000000;
slave_timing[3][27].info_i__max_slave__  = 0.027000000;
slave_timing[3][27].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][27].info_r__dsi_bus__    = 5.000;

slave_timing[3][27].t_rxd1[0][1] = 2824ns;
slave_timing[3][27].t_rxd1[1][0] = 3428ns;
slave_timing[3][27].t_rxd1[0][2] = 2179ns;
slave_timing[3][27].t_rxd1[2][0] = 3918ns;
slave_timing[3][27].t_rxd2[0][2] = 3189ns;
slave_timing[3][27].t_rxd2[2][0] = 2779ns;
slave_timing[3][27].t_rxd2[1][2] = 2277ns;
slave_timing[3][27].t_rxd2[2][1] = 4298ns;

slave_timing[3][28].info_corner          = 0;
slave_timing[3][28].info_temp__j__       = 25;
slave_timing[3][28].info_i__quite_rec__  = 0.003000000;
slave_timing[3][28].info_dtr__ib__       = 1;
slave_timing[3][28].info_i__offset_rec__ = -0.001000000;
slave_timing[3][28].info_i__max_slave__  = 0.021000000;
slave_timing[3][28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][28].info_r__dsi_bus__    = 5.000;

slave_timing[3][28].t_rxd1[0][1] = 3924ns;
slave_timing[3][28].t_rxd1[1][0] = 2671ns;
slave_timing[3][28].t_rxd1[0][2] = 2675ns;
slave_timing[3][28].t_rxd1[2][0] = 3413ns;
slave_timing[3][28].t_rxd2[0][2] = 4615ns;
slave_timing[3][28].t_rxd2[2][0] = 1983ns;
slave_timing[3][28].t_rxd2[1][2] = 4330ns;
slave_timing[3][28].t_rxd2[2][1] = 2518ns;

slave_timing[3][29].info_corner          = 0;
slave_timing[3][29].info_temp__j__       = 25;
slave_timing[3][29].info_i__quite_rec__  = 0.003000000;
slave_timing[3][29].info_dtr__ib__       = 1;
slave_timing[3][29].info_i__offset_rec__ = 0.001000000;
slave_timing[3][29].info_i__max_slave__  = 0.021000000;
slave_timing[3][29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][29].info_r__dsi_bus__    = 5.000;

slave_timing[3][29].t_rxd1[0][1] = 3290ns;
slave_timing[3][29].t_rxd1[1][0] = 3144ns;
slave_timing[3][29].t_rxd1[0][2] = 2435ns;
slave_timing[3][29].t_rxd1[2][0] = 3719ns;
slave_timing[3][29].t_rxd2[0][2] = 3975ns;
slave_timing[3][29].t_rxd2[2][0] = 2287ns;
slave_timing[3][29].t_rxd2[1][2] = 3508ns;
slave_timing[3][29].t_rxd2[2][1] = 2986ns;

slave_timing[3][30].info_corner          = 0;
slave_timing[3][30].info_temp__j__       = 25;
slave_timing[3][30].info_i__quite_rec__  = 0.003000000;
slave_timing[3][30].info_dtr__ib__       = 1;
slave_timing[3][30].info_i__offset_rec__ = -0.001000000;
slave_timing[3][30].info_i__max_slave__  = 0.027000000;
slave_timing[3][30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][30].info_r__dsi_bus__    = 5.000;

slave_timing[3][30].t_rxd1[0][1] = 3291ns;
slave_timing[3][30].t_rxd1[1][0] = 2974ns;
slave_timing[3][30].t_rxd1[0][2] = 2433ns;
slave_timing[3][30].t_rxd1[2][0] = 3604ns;
slave_timing[3][30].t_rxd2[0][2] = 3529ns;
slave_timing[3][30].t_rxd2[2][0] = 2509ns;
slave_timing[3][30].t_rxd2[1][2] = 2864ns;
slave_timing[3][30].t_rxd2[2][1] = 3441ns;

slave_timing[3][31].info_corner          = 0;
slave_timing[3][31].info_temp__j__       = 25;
slave_timing[3][31].info_i__quite_rec__  = 0.003000000;
slave_timing[3][31].info_dtr__ib__       = 1;
slave_timing[3][31].info_i__offset_rec__ = 0.001000000;
slave_timing[3][31].info_i__max_slave__  = 0.027000000;
slave_timing[3][31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][31].info_r__dsi_bus__    = 5.000;

slave_timing[3][31].t_rxd1[0][1] = 2940ns;
slave_timing[3][31].t_rxd1[1][0] = 3321ns;
slave_timing[3][31].t_rxd1[0][2] = 2251ns;
slave_timing[3][31].t_rxd1[2][0] = 3844ns;
slave_timing[3][31].t_rxd2[0][2] = 3328ns;
slave_timing[3][31].t_rxd2[2][0] = 2673ns;
slave_timing[3][31].t_rxd2[1][2] = 2547ns;
slave_timing[3][31].t_rxd2[2][1] = 3904ns;

slave_timing[3][32].info_corner          = 0;
slave_timing[3][32].info_temp__j__       = 25;
slave_timing[3][32].info_i__quite_rec__  = 0.000000000;
slave_timing[3][32].info_dtr__ib__       = -1;
slave_timing[3][32].info_i__offset_rec__ = -0.001000000;
slave_timing[3][32].info_i__max_slave__  = 0.021000000;
slave_timing[3][32].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][32].info_r__dsi_bus__    = 5.000;

slave_timing[3][32].t_rxd1[0][1] = 3540ns;
slave_timing[3][32].t_rxd1[1][0] = 2518ns;
slave_timing[3][32].t_rxd1[0][2] = 2425ns;
slave_timing[3][32].t_rxd1[2][0] = 3214ns;
slave_timing[3][32].t_rxd2[0][2] = 3942ns;
slave_timing[3][32].t_rxd2[2][0] = 1941ns;
slave_timing[3][32].t_rxd2[1][2] = 3571ns;
slave_timing[3][32].t_rxd2[2][1] = 2522ns;

slave_timing[3][33].info_corner          = 0;
slave_timing[3][33].info_temp__j__       = 25;
slave_timing[3][33].info_i__quite_rec__  = 0.000000000;
slave_timing[3][33].info_dtr__ib__       = -1;
slave_timing[3][33].info_i__offset_rec__ = 0.001000000;
slave_timing[3][33].info_i__max_slave__  = 0.021000000;
slave_timing[3][33].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][33].info_r__dsi_bus__    = 5.000;

slave_timing[3][33].t_rxd1[0][1] = 3016ns;
slave_timing[3][33].t_rxd1[1][0] = 2973ns;
slave_timing[3][33].t_rxd1[0][2] = 2191ns;
slave_timing[3][33].t_rxd1[2][0] = 3512ns;
slave_timing[3][33].t_rxd2[0][2] = 3522ns;
slave_timing[3][33].t_rxd2[2][0] = 2206ns;
slave_timing[3][33].t_rxd2[1][2] = 3037ns;
slave_timing[3][33].t_rxd2[2][1] = 2932ns;

slave_timing[3][34].info_corner          = 0;
slave_timing[3][34].info_temp__j__       = 25;
slave_timing[3][34].info_i__quite_rec__  = 0.000000000;
slave_timing[3][34].info_dtr__ib__       = -1;
slave_timing[3][34].info_i__offset_rec__ = -0.001000000;
slave_timing[3][34].info_i__max_slave__  = 0.027000000;
slave_timing[3][34].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][34].info_r__dsi_bus__    = 5.000;

slave_timing[3][34].t_rxd1[0][1] = 3028ns;
slave_timing[3][34].t_rxd1[1][0] = 2761ns;
slave_timing[3][34].t_rxd1[0][2] = 2220ns;
slave_timing[3][34].t_rxd1[2][0] = 3372ns;
slave_timing[3][34].t_rxd2[0][2] = 3193ns;
slave_timing[3][34].t_rxd2[2][0] = 2372ns;
slave_timing[3][34].t_rxd2[1][2] = 2505ns;
slave_timing[3][34].t_rxd2[2][1] = 3366ns;

slave_timing[3][35].info_corner          = 0;
slave_timing[3][35].info_temp__j__       = 25;
slave_timing[3][35].info_i__quite_rec__  = 0.000000000;
slave_timing[3][35].info_dtr__ib__       = -1;
slave_timing[3][35].info_i__offset_rec__ = 0.001000000;
slave_timing[3][35].info_i__max_slave__  = 0.027000000;
slave_timing[3][35].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][35].info_r__dsi_bus__    = 5.000;

slave_timing[3][35].t_rxd1[0][1] = 2665ns;
slave_timing[3][35].t_rxd1[1][0] = 3143ns;
slave_timing[3][35].t_rxd1[0][2] = 2018ns;
slave_timing[3][35].t_rxd1[2][0] = 3629ns;
slave_timing[3][35].t_rxd2[0][2] = 2991ns;
slave_timing[3][35].t_rxd2[2][0] = 2544ns;
slave_timing[3][35].t_rxd2[1][2] = 2144ns;
slave_timing[3][35].t_rxd2[2][1] = 3969ns;

slave_timing[3][36].info_corner          = 0;
slave_timing[3][36].info_temp__j__       = 25;
slave_timing[3][36].info_i__quite_rec__  = 0.000000000;
slave_timing[3][36].info_dtr__ib__       = 1;
slave_timing[3][36].info_i__offset_rec__ = -0.001000000;
slave_timing[3][36].info_i__max_slave__  = 0.021000000;
slave_timing[3][36].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][36].info_r__dsi_bus__    = 5.000;

slave_timing[3][36].t_rxd1[0][1] = 3806ns;
slave_timing[3][36].t_rxd1[1][0] = 2394ns;
slave_timing[3][36].t_rxd1[0][2] = 2503ns;
slave_timing[3][36].t_rxd1[2][0] = 3141ns;
slave_timing[3][36].t_rxd2[0][2] = 4509ns;
slave_timing[3][36].t_rxd2[2][0] = 1749ns;
slave_timing[3][36].t_rxd2[1][2] = 4296ns;
slave_timing[3][36].t_rxd2[2][1] = 2245ns;

slave_timing[3][37].info_corner          = 0;
slave_timing[3][37].info_temp__j__       = 25;
slave_timing[3][37].info_i__quite_rec__  = 0.000000000;
slave_timing[3][37].info_dtr__ib__       = 1;
slave_timing[3][37].info_i__offset_rec__ = 0.001000000;
slave_timing[3][37].info_i__max_slave__  = 0.021000000;
slave_timing[3][37].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][37].info_r__dsi_bus__    = 5.000;

slave_timing[3][37].t_rxd1[0][1] = 3149ns;
slave_timing[3][37].t_rxd1[1][0] = 2847ns;
slave_timing[3][37].t_rxd1[0][2] = 2276ns;
slave_timing[3][37].t_rxd1[2][0] = 3426ns;
slave_timing[3][37].t_rxd2[0][2] = 3790ns;
slave_timing[3][37].t_rxd2[2][0] = 2052ns;
slave_timing[3][37].t_rxd2[1][2] = 3368ns;
slave_timing[3][37].t_rxd2[2][1] = 2698ns;

slave_timing[3][38].info_corner          = 0;
slave_timing[3][38].info_temp__j__       = 25;
slave_timing[3][38].info_i__quite_rec__  = 0.000000000;
slave_timing[3][38].info_dtr__ib__       = 1;
slave_timing[3][38].info_i__offset_rec__ = -0.001000000;
slave_timing[3][38].info_i__max_slave__  = 0.027000000;
slave_timing[3][38].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][38].info_r__dsi_bus__    = 5.000;

slave_timing[3][38].t_rxd1[0][1] = 3130ns;
slave_timing[3][38].t_rxd1[1][0] = 2699ns;
slave_timing[3][38].t_rxd1[0][2] = 2267ns;
slave_timing[3][38].t_rxd1[2][0] = 3332ns;
slave_timing[3][38].t_rxd2[0][2] = 3328ns;
slave_timing[3][38].t_rxd2[2][0] = 2280ns;
slave_timing[3][38].t_rxd2[1][2] = 2708ns;
slave_timing[3][38].t_rxd2[2][1] = 3142ns;

slave_timing[3][39].info_corner          = 0;
slave_timing[3][39].info_temp__j__       = 25;
slave_timing[3][39].info_i__quite_rec__  = 0.000000000;
slave_timing[3][39].info_dtr__ib__       = 1;
slave_timing[3][39].info_i__offset_rec__ = 0.001000000;
slave_timing[3][39].info_i__max_slave__  = 0.027000000;
slave_timing[3][39].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][39].info_r__dsi_bus__    = 5.000;

slave_timing[3][39].t_rxd1[0][1] = 2752ns;
slave_timing[3][39].t_rxd1[1][0] = 3070ns;
slave_timing[3][39].t_rxd1[0][2] = 2074ns;
slave_timing[3][39].t_rxd1[2][0] = 3582ns;
slave_timing[3][39].t_rxd2[0][2] = 3111ns;
slave_timing[3][39].t_rxd2[2][0] = 2458ns;
slave_timing[3][39].t_rxd2[1][2] = 2366ns;
slave_timing[3][39].t_rxd2[2][1] = 3619ns;

slave_timing[3][40].info_corner          = 0;
slave_timing[3][40].info_temp__j__       = 25;
slave_timing[3][40].info_i__quite_rec__  = 0.000000000;
slave_timing[3][40].info_dtr__ib__       = -1;
slave_timing[3][40].info_i__offset_rec__ = -0.001000000;
slave_timing[3][40].info_i__max_slave__  = 0.021000000;
slave_timing[3][40].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][40].info_r__dsi_bus__    = 5.000;

slave_timing[3][40].t_rxd1[0][1] = 3777ns;
slave_timing[3][40].t_rxd1[1][0] = 2722ns;
slave_timing[3][40].t_rxd1[0][2] = 2652ns;
slave_timing[3][40].t_rxd1[2][0] = 3414ns;
slave_timing[3][40].t_rxd2[0][2] = 4264ns;
slave_timing[3][40].t_rxd2[2][0] = 2104ns;
slave_timing[3][40].t_rxd2[1][2] = 3815ns;
slave_timing[3][40].t_rxd2[2][1] = 2730ns;

slave_timing[3][41].info_corner          = 0;
slave_timing[3][41].info_temp__j__       = 25;
slave_timing[3][41].info_i__quite_rec__  = 0.000000000;
slave_timing[3][41].info_dtr__ib__       = -1;
slave_timing[3][41].info_i__offset_rec__ = 0.001000000;
slave_timing[3][41].info_i__max_slave__  = 0.021000000;
slave_timing[3][41].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][41].info_r__dsi_bus__    = 5.000;

slave_timing[3][41].t_rxd1[0][1] = 3194ns;
slave_timing[3][41].t_rxd1[1][0] = 3196ns;
slave_timing[3][41].t_rxd1[0][2] = 2388ns;
slave_timing[3][41].t_rxd1[2][0] = 3756ns;
slave_timing[3][41].t_rxd2[0][2] = 3766ns;
slave_timing[3][41].t_rxd2[2][0] = 2402ns;
slave_timing[3][41].t_rxd2[1][2] = 3217ns;
slave_timing[3][41].t_rxd2[2][1] = 3204ns;

slave_timing[3][42].info_corner          = 0;
slave_timing[3][42].info_temp__j__       = 25;
slave_timing[3][42].info_i__quite_rec__  = 0.000000000;
slave_timing[3][42].info_dtr__ib__       = -1;
slave_timing[3][42].info_i__offset_rec__ = -0.001000000;
slave_timing[3][42].info_i__max_slave__  = 0.027000000;
slave_timing[3][42].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][42].info_r__dsi_bus__    = 5.000;

slave_timing[3][42].t_rxd1[0][1] = 3257ns;
slave_timing[3][42].t_rxd1[1][0] = 2980ns;
slave_timing[3][42].t_rxd1[0][2] = 2414ns;
slave_timing[3][42].t_rxd1[2][0] = 3609ns;
slave_timing[3][42].t_rxd2[0][2] = 3428ns;
slave_timing[3][42].t_rxd2[2][0] = 2572ns;
slave_timing[3][42].t_rxd2[1][2] = 2713ns;
slave_timing[3][42].t_rxd2[2][1] = 3605ns;

slave_timing[3][43].info_corner          = 0;
slave_timing[3][43].info_temp__j__       = 25;
slave_timing[3][43].info_i__quite_rec__  = 0.000000000;
slave_timing[3][43].info_dtr__ib__       = -1;
slave_timing[3][43].info_i__offset_rec__ = 0.001000000;
slave_timing[3][43].info_i__max_slave__  = 0.027000000;
slave_timing[3][43].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][43].info_r__dsi_bus__    = 5.000;

slave_timing[3][43].t_rxd1[0][1] = 2879ns;
slave_timing[3][43].t_rxd1[1][0] = 3371ns;
slave_timing[3][43].t_rxd1[0][2] = 2210ns;
slave_timing[3][43].t_rxd1[2][0] = 3878ns;
slave_timing[3][43].t_rxd2[0][2] = 3214ns;
slave_timing[3][43].t_rxd2[2][0] = 2754ns;
slave_timing[3][43].t_rxd2[1][2] = 2340ns;
slave_timing[3][43].t_rxd2[2][1] = 4243ns;

slave_timing[3][44].info_corner          = 0;
slave_timing[3][44].info_temp__j__       = 25;
slave_timing[3][44].info_i__quite_rec__  = 0.000000000;
slave_timing[3][44].info_dtr__ib__       = 1;
slave_timing[3][44].info_i__offset_rec__ = -0.001000000;
slave_timing[3][44].info_i__max_slave__  = 0.021000000;
slave_timing[3][44].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][44].info_r__dsi_bus__    = 5.000;

slave_timing[3][44].t_rxd1[0][1] = 3979ns;
slave_timing[3][44].t_rxd1[1][0] = 2645ns;
slave_timing[3][44].t_rxd1[0][2] = 2713ns;
slave_timing[3][44].t_rxd1[2][0] = 3369ns;
slave_timing[3][44].t_rxd2[0][2] = 4820ns;
slave_timing[3][44].t_rxd2[2][0] = 1936ns;
slave_timing[3][44].t_rxd2[1][2] = 4400ns;
slave_timing[3][44].t_rxd2[2][1] = 2488ns;

slave_timing[3][45].info_corner          = 0;
slave_timing[3][45].info_temp__j__       = 25;
slave_timing[3][45].info_i__quite_rec__  = 0.000000000;
slave_timing[3][45].info_dtr__ib__       = 1;
slave_timing[3][45].info_i__offset_rec__ = 0.001000000;
slave_timing[3][45].info_i__max_slave__  = 0.021000000;
slave_timing[3][45].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][45].info_r__dsi_bus__    = 5.000;

slave_timing[3][45].t_rxd1[0][1] = 3323ns;
slave_timing[3][45].t_rxd1[1][0] = 3116ns;
slave_timing[3][45].t_rxd1[0][2] = 2450ns;
slave_timing[3][45].t_rxd1[2][0] = 3700ns;
slave_timing[3][45].t_rxd2[0][2] = 4001ns;
slave_timing[3][45].t_rxd2[2][0] = 2271ns;
slave_timing[3][45].t_rxd2[1][2] = 3544ns;
slave_timing[3][45].t_rxd2[2][1] = 2956ns;

slave_timing[3][46].info_corner          = 0;
slave_timing[3][46].info_temp__j__       = 25;
slave_timing[3][46].info_i__quite_rec__  = 0.000000000;
slave_timing[3][46].info_dtr__ib__       = 1;
slave_timing[3][46].info_i__offset_rec__ = -0.001000000;
slave_timing[3][46].info_i__max_slave__  = 0.027000000;
slave_timing[3][46].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][46].info_r__dsi_bus__    = 5.000;

slave_timing[3][46].t_rxd1[0][1] = 3361ns;
slave_timing[3][46].t_rxd1[1][0] = 2916ns;
slave_timing[3][46].t_rxd1[0][2] = 2464ns;
slave_timing[3][46].t_rxd1[2][0] = 3565ns;
slave_timing[3][46].t_rxd2[0][2] = 3566ns;
slave_timing[3][46].t_rxd2[2][0] = 2476ns;
slave_timing[3][46].t_rxd2[1][2] = 2928ns;
slave_timing[3][46].t_rxd2[2][1] = 3369ns;

slave_timing[3][47].info_corner          = 0;
slave_timing[3][47].info_temp__j__       = 25;
slave_timing[3][47].info_i__quite_rec__  = 0.000000000;
slave_timing[3][47].info_dtr__ib__       = 1;
slave_timing[3][47].info_i__offset_rec__ = 0.001000000;
slave_timing[3][47].info_i__max_slave__  = 0.027000000;
slave_timing[3][47].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][47].info_r__dsi_bus__    = 5.000;

slave_timing[3][47].t_rxd1[0][1] = 2969ns;
slave_timing[3][47].t_rxd1[1][0] = 3299ns;
slave_timing[3][47].t_rxd1[0][2] = 2264ns;
slave_timing[3][47].t_rxd1[2][0] = 3829ns;
slave_timing[3][47].t_rxd2[0][2] = 3342ns;
slave_timing[3][47].t_rxd2[2][0] = 2662ns;
slave_timing[3][47].t_rxd2[1][2] = 2569ns;
slave_timing[3][47].t_rxd2[2][1] = 3872ns;

slave_timing[3][48].info_corner          = 0;
slave_timing[3][48].info_temp__j__       = 25;
slave_timing[3][48].info_i__quite_rec__  = 0.040000000;
slave_timing[3][48].info_dtr__ib__       = -1;
slave_timing[3][48].info_i__offset_rec__ = -0.001000000;
slave_timing[3][48].info_i__max_slave__  = 0.021000000;
slave_timing[3][48].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][48].info_r__dsi_bus__    = 5.000;

slave_timing[3][48].t_rxd1[0][1] = 3331ns;
slave_timing[3][48].t_rxd1[1][0] = 2659ns;
slave_timing[3][48].t_rxd1[0][2] = 2353ns;
slave_timing[3][48].t_rxd1[2][0] = 3306ns;
slave_timing[3][48].t_rxd2[0][2] = 3788ns;
slave_timing[3][48].t_rxd2[2][0] = 2031ns;
slave_timing[3][48].t_rxd2[1][2] = 3366ns;
slave_timing[3][48].t_rxd2[2][1] = 2657ns;

slave_timing[3][49].info_corner          = 0;
slave_timing[3][49].info_temp__j__       = 25;
slave_timing[3][49].info_i__quite_rec__  = 0.040000000;
slave_timing[3][49].info_dtr__ib__       = -1;
slave_timing[3][49].info_i__offset_rec__ = 0.001000000;
slave_timing[3][49].info_i__max_slave__  = 0.021000000;
slave_timing[3][49].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][49].info_r__dsi_bus__    = 5.000;

slave_timing[3][49].t_rxd1[0][1] = 2820ns;
slave_timing[3][49].t_rxd1[1][0] = 3129ns;
slave_timing[3][49].t_rxd1[0][2] = 2113ns;
slave_timing[3][49].t_rxd1[2][0] = 3629ns;
slave_timing[3][49].t_rxd2[0][2] = 3413ns;
slave_timing[3][49].t_rxd2[2][0] = 2281ns;
slave_timing[3][49].t_rxd2[1][2] = 2841ns;
slave_timing[3][49].t_rxd2[2][1] = 3133ns;

slave_timing[3][50].info_corner          = 0;
slave_timing[3][50].info_temp__j__       = 25;
slave_timing[3][50].info_i__quite_rec__  = 0.040000000;
slave_timing[3][50].info_dtr__ib__       = -1;
slave_timing[3][50].info_i__offset_rec__ = -0.001000000;
slave_timing[3][50].info_i__max_slave__  = 0.027000000;
slave_timing[3][50].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][50].info_r__dsi_bus__    = 5.000;

slave_timing[3][50].t_rxd1[0][1] = 2942ns;
slave_timing[3][50].t_rxd1[1][0] = 2845ns;
slave_timing[3][50].t_rxd1[0][2] = 2177ns;
slave_timing[3][50].t_rxd1[2][0] = 3425ns;
slave_timing[3][50].t_rxd2[0][2] = 3145ns;
slave_timing[3][50].t_rxd2[2][0] = 2408ns;
slave_timing[3][50].t_rxd2[1][2] = 2431ns;
slave_timing[3][50].t_rxd2[2][1] = 3468ns;

slave_timing[3][51].info_corner          = 0;
slave_timing[3][51].info_temp__j__       = 25;
slave_timing[3][51].info_i__quite_rec__  = 0.040000000;
slave_timing[3][51].info_dtr__ib__       = -1;
slave_timing[3][51].info_i__offset_rec__ = 0.001000000;
slave_timing[3][51].info_i__max_slave__  = 0.027000000;
slave_timing[3][51].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][51].info_r__dsi_bus__    = 5.000;

slave_timing[3][51].t_rxd1[0][1] = 2622ns;
slave_timing[3][51].t_rxd1[1][0] = 3195ns;
slave_timing[3][51].t_rxd1[0][2] = 1991ns;
slave_timing[3][51].t_rxd1[2][0] = 3674ns;
slave_timing[3][51].t_rxd2[0][2] = 2966ns;
slave_timing[3][51].t_rxd2[2][0] = 2565ns;
slave_timing[3][51].t_rxd2[1][2] = 2094ns;
slave_timing[3][51].t_rxd2[2][1] = 4090ns;

slave_timing[3][52].info_corner          = 0;
slave_timing[3][52].info_temp__j__       = 25;
slave_timing[3][52].info_i__quite_rec__  = 0.040000000;
slave_timing[3][52].info_dtr__ib__       = 1;
slave_timing[3][52].info_i__offset_rec__ = -0.001000000;
slave_timing[3][52].info_i__max_slave__  = 0.021000000;
slave_timing[3][52].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][52].info_r__dsi_bus__    = 5.000;

slave_timing[3][52].t_rxd1[0][1] = 3745ns;
slave_timing[3][52].t_rxd1[1][0] = 2427ns;
slave_timing[3][52].t_rxd1[0][2] = 2487ns;
slave_timing[3][52].t_rxd1[2][0] = 3162ns;
slave_timing[3][52].t_rxd2[0][2] = 4414ns;
slave_timing[3][52].t_rxd2[2][0] = 1772ns;
slave_timing[3][52].t_rxd2[1][2] = 4176ns;
slave_timing[3][52].t_rxd2[2][1] = 2280ns;

slave_timing[3][53].info_corner          = 0;
slave_timing[3][53].info_temp__j__       = 25;
slave_timing[3][53].info_i__quite_rec__  = 0.040000000;
slave_timing[3][53].info_dtr__ib__       = 1;
slave_timing[3][53].info_i__offset_rec__ = 0.001000000;
slave_timing[3][53].info_i__max_slave__  = 0.021000000;
slave_timing[3][53].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][53].info_r__dsi_bus__    = 5.000;

slave_timing[3][53].t_rxd1[0][1] = 3108ns;
slave_timing[3][53].t_rxd1[1][0] = 2877ns;
slave_timing[3][53].t_rxd1[0][2] = 2255ns;
slave_timing[3][53].t_rxd1[2][0] = 3450ns;
slave_timing[3][53].t_rxd2[0][2] = 3755ns;
slave_timing[3][53].t_rxd2[2][0] = 2070ns;
slave_timing[3][53].t_rxd2[1][2] = 3320ns;
slave_timing[3][53].t_rxd2[2][1] = 2682ns;

slave_timing[3][54].info_corner          = 0;
slave_timing[3][54].info_temp__j__       = 25;
slave_timing[3][54].info_i__quite_rec__  = 0.040000000;
slave_timing[3][54].info_dtr__ib__       = 1;
slave_timing[3][54].info_i__offset_rec__ = -0.001000000;
slave_timing[3][54].info_i__max_slave__  = 0.027000000;
slave_timing[3][54].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][54].info_r__dsi_bus__    = 5.000;

slave_timing[3][54].t_rxd1[0][1] = 3141ns;
slave_timing[3][54].t_rxd1[1][0] = 2690ns;
slave_timing[3][54].t_rxd1[0][2] = 2272ns;
slave_timing[3][54].t_rxd1[2][0] = 3325ns;
slave_timing[3][54].t_rxd2[0][2] = 3334ns;
slave_timing[3][54].t_rxd2[2][0] = 2275ns;
slave_timing[3][54].t_rxd2[1][2] = 2722ns;
slave_timing[3][54].t_rxd2[2][1] = 3127ns;

slave_timing[3][55].info_corner          = 0;
slave_timing[3][55].info_temp__j__       = 25;
slave_timing[3][55].info_i__quite_rec__  = 0.040000000;
slave_timing[3][55].info_dtr__ib__       = 1;
slave_timing[3][55].info_i__offset_rec__ = 0.001000000;
slave_timing[3][55].info_i__max_slave__  = 0.027000000;
slave_timing[3][55].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][55].info_r__dsi_bus__    = 5.000;

slave_timing[3][55].t_rxd1[0][1] = 2761ns;
slave_timing[3][55].t_rxd1[1][0] = 3058ns;
slave_timing[3][55].t_rxd1[0][2] = 2079ns;
slave_timing[3][55].t_rxd1[2][0] = 3572ns;
slave_timing[3][55].t_rxd2[0][2] = 3115ns;
slave_timing[3][55].t_rxd2[2][0] = 2450ns;
slave_timing[3][55].t_rxd2[1][2] = 2376ns;
slave_timing[3][55].t_rxd2[2][1] = 3608ns;

slave_timing[3][56].info_corner          = 0;
slave_timing[3][56].info_temp__j__       = 25;
slave_timing[3][56].info_i__quite_rec__  = 0.040000000;
slave_timing[3][56].info_dtr__ib__       = -1;
slave_timing[3][56].info_i__offset_rec__ = -0.001000000;
slave_timing[3][56].info_i__max_slave__  = 0.021000000;
slave_timing[3][56].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][56].info_r__dsi_bus__    = 5.000;

slave_timing[3][56].t_rxd1[0][1] = 3569ns;
slave_timing[3][56].t_rxd1[1][0] = 2868ns;
slave_timing[3][56].t_rxd1[0][2] = 2556ns;
slave_timing[3][56].t_rxd1[2][0] = 3538ns;
slave_timing[3][56].t_rxd2[0][2] = 4044ns;
slave_timing[3][56].t_rxd2[2][0] = 2220ns;
slave_timing[3][56].t_rxd2[1][2] = 3603ns;
slave_timing[3][56].t_rxd2[2][1] = 2873ns;

slave_timing[3][57].info_corner          = 0;
slave_timing[3][57].info_temp__j__       = 25;
slave_timing[3][57].info_i__quite_rec__  = 0.040000000;
slave_timing[3][57].info_dtr__ib__       = -1;
slave_timing[3][57].info_i__offset_rec__ = 0.001000000;
slave_timing[3][57].info_i__max_slave__  = 0.021000000;
slave_timing[3][57].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][57].info_r__dsi_bus__    = 5.000;

slave_timing[3][57].t_rxd1[0][1] = 3082ns;
slave_timing[3][57].t_rxd1[1][0] = 3314ns;
slave_timing[3][57].t_rxd1[0][2] = 2305ns;
slave_timing[3][57].t_rxd1[2][0] = 3841ns;
slave_timing[3][57].t_rxd2[0][2] = 3657ns;
slave_timing[3][57].t_rxd2[2][0] = 2454ns;
slave_timing[3][57].t_rxd2[1][2] = 3109ns;
slave_timing[3][57].t_rxd2[2][1] = 3303ns;

slave_timing[3][58].info_corner          = 0;
slave_timing[3][58].info_temp__j__       = 25;
slave_timing[3][58].info_i__quite_rec__  = 0.040000000;
slave_timing[3][58].info_dtr__ib__       = -1;
slave_timing[3][58].info_i__offset_rec__ = -0.001000000;
slave_timing[3][58].info_i__max_slave__  = 0.027000000;
slave_timing[3][58].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][58].info_r__dsi_bus__    = 5.000;

slave_timing[3][58].t_rxd1[0][1] = 3168ns;
slave_timing[3][58].t_rxd1[1][0] = 3069ns;
slave_timing[3][58].t_rxd1[0][2] = 2374ns;
slave_timing[3][58].t_rxd1[2][0] = 3666ns;
slave_timing[3][58].t_rxd2[0][2] = 3381ns;
slave_timing[3][58].t_rxd2[2][0] = 2611ns;
slave_timing[3][58].t_rxd2[1][2] = 2633ns;
slave_timing[3][58].t_rxd2[2][1] = 3714ns;

slave_timing[3][59].info_corner          = 0;
slave_timing[3][59].info_temp__j__       = 25;
slave_timing[3][59].info_i__quite_rec__  = 0.040000000;
slave_timing[3][59].info_dtr__ib__       = -1;
slave_timing[3][59].info_i__offset_rec__ = 0.001000000;
slave_timing[3][59].info_i__max_slave__  = 0.027000000;
slave_timing[3][59].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][59].info_r__dsi_bus__    = 5.000;

slave_timing[3][59].t_rxd1[0][1] = 2829ns;
slave_timing[3][59].t_rxd1[1][0] = 3429ns;
slave_timing[3][59].t_rxd1[0][2] = 2183ns;
slave_timing[3][59].t_rxd1[2][0] = 3924ns;
slave_timing[3][59].t_rxd2[0][2] = 3191ns;
slave_timing[3][59].t_rxd2[2][0] = 2776ns;
slave_timing[3][59].t_rxd2[1][2] = 2283ns;
slave_timing[3][59].t_rxd2[2][1] = 4379ns;

slave_timing[3][60].info_corner          = 0;
slave_timing[3][60].info_temp__j__       = 25;
slave_timing[3][60].info_i__quite_rec__  = 0.040000000;
slave_timing[3][60].info_dtr__ib__       = 1;
slave_timing[3][60].info_i__offset_rec__ = -0.001000000;
slave_timing[3][60].info_i__max_slave__  = 0.021000000;
slave_timing[3][60].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][60].info_r__dsi_bus__    = 5.000;

slave_timing[3][60].t_rxd1[0][1] = 4003ns;
slave_timing[3][60].t_rxd1[1][0] = 2631ns;
slave_timing[3][60].t_rxd1[0][2] = 2694ns;
slave_timing[3][60].t_rxd1[2][0] = 3390ns;
slave_timing[3][60].t_rxd2[0][2] = 4725ns;
slave_timing[3][60].t_rxd2[2][0] = 1961ns;
slave_timing[3][60].t_rxd2[1][2] = 4446ns;
slave_timing[3][60].t_rxd2[2][1] = 2480ns;

slave_timing[3][61].info_corner          = 0;
slave_timing[3][61].info_temp__j__       = 25;
slave_timing[3][61].info_i__quite_rec__  = 0.040000000;
slave_timing[3][61].info_dtr__ib__       = 1;
slave_timing[3][61].info_i__offset_rec__ = 0.001000000;
slave_timing[3][61].info_i__max_slave__  = 0.021000000;
slave_timing[3][61].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][61].info_r__dsi_bus__    = 5.000;

slave_timing[3][61].t_rxd1[0][1] = 3335ns;
slave_timing[3][61].t_rxd1[1][0] = 3099ns;
slave_timing[3][61].t_rxd1[0][2] = 2456ns;
slave_timing[3][61].t_rxd1[2][0] = 3691ns;
slave_timing[3][61].t_rxd2[0][2] = 4015ns;
slave_timing[3][61].t_rxd2[2][0] = 2265ns;
slave_timing[3][61].t_rxd2[1][2] = 3561ns;
slave_timing[3][61].t_rxd2[2][1] = 2945ns;

slave_timing[3][62].info_corner          = 0;
slave_timing[3][62].info_temp__j__       = 25;
slave_timing[3][62].info_i__quite_rec__  = 0.040000000;
slave_timing[3][62].info_dtr__ib__       = 1;
slave_timing[3][62].info_i__offset_rec__ = -0.001000000;
slave_timing[3][62].info_i__max_slave__  = 0.027000000;
slave_timing[3][62].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][62].info_r__dsi_bus__    = 5.000;

slave_timing[3][62].t_rxd1[0][1] = 3373ns;
slave_timing[3][62].t_rxd1[1][0] = 2903ns;
slave_timing[3][62].t_rxd1[0][2] = 2478ns;
slave_timing[3][62].t_rxd1[2][0] = 3560ns;
slave_timing[3][62].t_rxd2[0][2] = 3580ns;
slave_timing[3][62].t_rxd2[2][0] = 2471ns;
slave_timing[3][62].t_rxd2[1][2] = 2940ns;
slave_timing[3][62].t_rxd2[2][1] = 3360ns;

slave_timing[3][63].info_corner          = 0;
slave_timing[3][63].info_temp__j__       = 25;
slave_timing[3][63].info_i__quite_rec__  = 0.040000000;
slave_timing[3][63].info_dtr__ib__       = 1;
slave_timing[3][63].info_i__offset_rec__ = 0.001000000;
slave_timing[3][63].info_i__max_slave__  = 0.027000000;
slave_timing[3][63].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][63].info_r__dsi_bus__    = 5.000;

slave_timing[3][63].t_rxd1[0][1] = 2981ns;
slave_timing[3][63].t_rxd1[1][0] = 3286ns;
slave_timing[3][63].t_rxd1[0][2] = 2273ns;
slave_timing[3][63].t_rxd1[2][0] = 3820ns;
slave_timing[3][63].t_rxd2[0][2] = 3347ns;
slave_timing[3][63].t_rxd2[2][0] = 2658ns;
slave_timing[3][63].t_rxd2[1][2] = 2577ns;
slave_timing[3][63].t_rxd2[2][1] = 3850ns;


slave_timing[2][64+0].info_corner          = 3;
slave_timing[2][64+0].info_temp__j__       = 125;
slave_timing[2][64+0].info_i__quite_rec__  = 0.006000000;
slave_timing[2][64+0].info_dtr__ib__       = -1;
slave_timing[2][64+0].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+0].info_i__max_slave__  = 0.023000000;
slave_timing[2][64+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][64+0].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+0].t_rxd1[0][1] = 2196ns;
slave_timing[2][64+0].t_rxd1[1][0] = 2166ns;
slave_timing[2][64+0].t_rxd1[0][2] = 1641ns;
slave_timing[2][64+0].t_rxd1[2][0] = 2644ns;
slave_timing[2][64+0].t_rxd2[0][2] = 2622ns;
slave_timing[2][64+0].t_rxd2[2][0] = 1659ns;
slave_timing[2][64+0].t_rxd2[1][2] = 2204ns;
slave_timing[2][64+0].t_rxd2[2][1] = 2177ns;

slave_timing[2][64+1].info_corner          = 3;
slave_timing[2][64+1].info_temp__j__       = 125;
slave_timing[2][64+1].info_i__quite_rec__  = 0.006000000;
slave_timing[2][64+1].info_dtr__ib__       = -1;
slave_timing[2][64+1].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+1].info_i__max_slave__  = 0.025000000;
slave_timing[2][64+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][64+1].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+1].t_rxd1[0][1] = 2102ns;
slave_timing[2][64+1].t_rxd1[1][0] = 2241ns;
slave_timing[2][64+1].t_rxd1[0][2] = 1610ns;
slave_timing[2][64+1].t_rxd1[2][0] = 2689ns;
slave_timing[2][64+1].t_rxd2[0][2] = 2489ns;
slave_timing[2][64+1].t_rxd2[2][0] = 1773ns;
slave_timing[2][64+1].t_rxd2[1][2] = 1961ns;
slave_timing[2][64+1].t_rxd2[2][1] = 2403ns;

slave_timing[2][64+2].info_corner          = 3;
slave_timing[2][64+2].info_temp__j__       = 125;
slave_timing[2][64+2].info_i__quite_rec__  = 0.006000000;
slave_timing[2][64+2].info_dtr__ib__       = 1;
slave_timing[2][64+2].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+2].info_i__max_slave__  = 0.023000000;
slave_timing[2][64+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][64+2].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+2].t_rxd1[0][1] = 2233ns;
slave_timing[2][64+2].t_rxd1[1][0] = 2110ns;
slave_timing[2][64+2].t_rxd1[0][2] = 1674ns;
slave_timing[2][64+2].t_rxd1[2][0] = 2584ns;
slave_timing[2][64+2].t_rxd2[0][2] = 2756ns;
slave_timing[2][64+2].t_rxd2[2][0] = 1538ns;
slave_timing[2][64+2].t_rxd2[1][2] = 2376ns;
slave_timing[2][64+2].t_rxd2[2][1] = 1983ns;

slave_timing[2][64+3].info_corner          = 3;
slave_timing[2][64+3].info_temp__j__       = 125;
slave_timing[2][64+3].info_i__quite_rec__  = 0.006000000;
slave_timing[2][64+3].info_dtr__ib__       = 1;
slave_timing[2][64+3].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+3].info_i__max_slave__  = 0.025000000;
slave_timing[2][64+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][64+3].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+3].t_rxd1[0][1] = 2145ns;
slave_timing[2][64+3].t_rxd1[1][0] = 2169ns;
slave_timing[2][64+3].t_rxd1[0][2] = 1623ns;
slave_timing[2][64+3].t_rxd1[2][0] = 2626ns;
slave_timing[2][64+3].t_rxd2[0][2] = 2579ns;
slave_timing[2][64+3].t_rxd2[2][0] = 1678ns;
slave_timing[2][64+3].t_rxd2[1][2] = 2123ns;
slave_timing[2][64+3].t_rxd2[2][1] = 2214ns;

slave_timing[2][64+4].info_corner          = 3;
slave_timing[2][64+4].info_temp__j__       = 125;
slave_timing[2][64+4].info_i__quite_rec__  = 0.006000000;
slave_timing[2][64+4].info_dtr__ib__       = -1;
slave_timing[2][64+4].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+4].info_i__max_slave__  = 0.023000000;
slave_timing[2][64+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][64+4].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+4].t_rxd1[0][1] = 2392ns;
slave_timing[2][64+4].t_rxd1[1][0] = 2327ns;
slave_timing[2][64+4].t_rxd1[0][2] = 1825ns;
slave_timing[2][64+4].t_rxd1[2][0] = 2788ns;
slave_timing[2][64+4].t_rxd2[0][2] = 2675ns;
slave_timing[2][64+4].t_rxd2[2][0] = 1694ns;
slave_timing[2][64+4].t_rxd2[1][2] = 2230ns;
slave_timing[2][64+4].t_rxd2[2][1] = 2207ns;

slave_timing[2][64+5].info_corner          = 3;
slave_timing[2][64+5].info_temp__j__       = 125;
slave_timing[2][64+5].info_i__quite_rec__  = 0.006000000;
slave_timing[2][64+5].info_dtr__ib__       = -1;
slave_timing[2][64+5].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+5].info_i__max_slave__  = 0.025000000;
slave_timing[2][64+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][64+5].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+5].t_rxd1[0][1] = 2308ns;
slave_timing[2][64+5].t_rxd1[1][0] = 2393ns;
slave_timing[2][64+5].t_rxd1[0][2] = 1772ns;
slave_timing[2][64+5].t_rxd1[2][0] = 2830ns;
slave_timing[2][64+5].t_rxd2[0][2] = 2530ns;
slave_timing[2][64+5].t_rxd2[2][0] = 1805ns;
slave_timing[2][64+5].t_rxd2[1][2] = 2001ns;
slave_timing[2][64+5].t_rxd2[2][1] = 2430ns;

slave_timing[2][64+6].info_corner          = 3;
slave_timing[2][64+6].info_temp__j__       = 125;
slave_timing[2][64+6].info_i__quite_rec__  = 0.006000000;
slave_timing[2][64+6].info_dtr__ib__       = 1;
slave_timing[2][64+6].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+6].info_i__max_slave__  = 0.023000000;
slave_timing[2][64+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][64+6].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+6].t_rxd1[0][1] = 2414ns;
slave_timing[2][64+6].t_rxd1[1][0] = 2245ns;
slave_timing[2][64+6].t_rxd1[0][2] = 1832ns;
slave_timing[2][64+6].t_rxd1[2][0] = 2722ns;
slave_timing[2][64+6].t_rxd2[0][2] = 2792ns;
slave_timing[2][64+6].t_rxd2[2][0] = 1573ns;
slave_timing[2][64+6].t_rxd2[1][2] = 2403ns;
slave_timing[2][64+6].t_rxd2[2][1] = 2017ns;

slave_timing[2][64+7].info_corner          = 3;
slave_timing[2][64+7].info_temp__j__       = 125;
slave_timing[2][64+7].info_i__quite_rec__  = 0.006000000;
slave_timing[2][64+7].info_dtr__ib__       = 1;
slave_timing[2][64+7].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+7].info_i__max_slave__  = 0.025000000;
slave_timing[2][64+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][64+7].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+7].t_rxd1[0][1] = 2327ns;
slave_timing[2][64+7].t_rxd1[1][0] = 2316ns;
slave_timing[2][64+7].t_rxd1[0][2] = 1781ns;
slave_timing[2][64+7].t_rxd1[2][0] = 2765ns;
slave_timing[2][64+7].t_rxd2[0][2] = 2617ns;
slave_timing[2][64+7].t_rxd2[2][0] = 1704ns;
slave_timing[2][64+7].t_rxd2[1][2] = 2142ns;
slave_timing[2][64+7].t_rxd2[2][1] = 2210ns;

slave_timing[2][64+8].info_corner          = 3;
slave_timing[2][64+8].info_temp__j__       = 125;
slave_timing[2][64+8].info_i__quite_rec__  = 0.003000000;
slave_timing[2][64+8].info_dtr__ib__       = -1;
slave_timing[2][64+8].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+8].info_i__max_slave__  = 0.023000000;
slave_timing[2][64+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][64+8].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+8].t_rxd1[0][1] = 2134ns;
slave_timing[2][64+8].t_rxd1[1][0] = 2164ns;
slave_timing[2][64+8].t_rxd1[0][2] = 1617ns;
slave_timing[2][64+8].t_rxd1[2][0] = 2618ns;
slave_timing[2][64+8].t_rxd2[0][2] = 2598ns;
slave_timing[2][64+8].t_rxd2[2][0] = 1647ns;
slave_timing[2][64+8].t_rxd2[1][2] = 2145ns;
slave_timing[2][64+8].t_rxd2[2][1] = 2159ns;

slave_timing[2][64+9].info_corner          = 3;
slave_timing[2][64+9].info_temp__j__       = 125;
slave_timing[2][64+9].info_i__quite_rec__  = 0.003000000;
slave_timing[2][64+9].info_dtr__ib__       = -1;
slave_timing[2][64+9].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+9].info_i__max_slave__  = 0.025000000;
slave_timing[2][64+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][64+9].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+9].t_rxd1[0][1] = 2057ns;
slave_timing[2][64+9].t_rxd1[1][0] = 2231ns;
slave_timing[2][64+9].t_rxd1[0][2] = 1572ns;
slave_timing[2][64+9].t_rxd1[2][0] = 2662ns;
slave_timing[2][64+9].t_rxd2[0][2] = 2448ns;
slave_timing[2][64+9].t_rxd2[2][0] = 1758ns;
slave_timing[2][64+9].t_rxd2[1][2] = 1922ns;
slave_timing[2][64+9].t_rxd2[2][1] = 2387ns;

slave_timing[2][64+10].info_corner          = 3;
slave_timing[2][64+10].info_temp__j__       = 125;
slave_timing[2][64+10].info_i__quite_rec__  = 0.003000000;
slave_timing[2][64+10].info_dtr__ib__       = 1;
slave_timing[2][64+10].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+10].info_i__max_slave__  = 0.023000000;
slave_timing[2][64+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][64+10].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+10].t_rxd1[0][1] = 2209ns;
slave_timing[2][64+10].t_rxd1[1][0] = 2061ns;
slave_timing[2][64+10].t_rxd1[0][2] = 1650ns;
slave_timing[2][64+10].t_rxd1[2][0] = 2536ns;
slave_timing[2][64+10].t_rxd2[0][2] = 2734ns;
slave_timing[2][64+10].t_rxd2[2][0] = 1514ns;
slave_timing[2][64+10].t_rxd2[1][2] = 2373ns;
slave_timing[2][64+10].t_rxd2[2][1] = 1945ns;

slave_timing[2][64+11].info_corner          = 3;
slave_timing[2][64+11].info_temp__j__       = 125;
slave_timing[2][64+11].info_i__quite_rec__  = 0.003000000;
slave_timing[2][64+11].info_dtr__ib__       = 1;
slave_timing[2][64+11].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+11].info_i__max_slave__  = 0.025000000;
slave_timing[2][64+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][64+11].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+11].t_rxd1[0][1] = 2111ns;
slave_timing[2][64+11].t_rxd1[1][0] = 2126ns;
slave_timing[2][64+11].t_rxd1[0][2] = 1597ns;
slave_timing[2][64+11].t_rxd1[2][0] = 2578ns;
slave_timing[2][64+11].t_rxd2[0][2] = 2558ns;
slave_timing[2][64+11].t_rxd2[2][0] = 1642ns;
slave_timing[2][64+11].t_rxd2[1][2] = 2103ns;
slave_timing[2][64+11].t_rxd2[2][1] = 2171ns;

slave_timing[2][64+12].info_corner          = 3;
slave_timing[2][64+12].info_temp__j__       = 125;
slave_timing[2][64+12].info_i__quite_rec__  = 0.003000000;
slave_timing[2][64+12].info_dtr__ib__       = -1;
slave_timing[2][64+12].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+12].info_i__max_slave__  = 0.023000000;
slave_timing[2][64+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][64+12].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+12].t_rxd1[0][1] = 2350ns;
slave_timing[2][64+12].t_rxd1[1][0] = 2323ns;
slave_timing[2][64+12].t_rxd1[0][2] = 1799ns;
slave_timing[2][64+12].t_rxd1[2][0] = 2770ns;
slave_timing[2][64+12].t_rxd2[0][2] = 2633ns;
slave_timing[2][64+12].t_rxd2[2][0] = 1675ns;
slave_timing[2][64+12].t_rxd2[1][2] = 2212ns;
slave_timing[2][64+12].t_rxd2[2][1] = 2133ns;

slave_timing[2][64+13].info_corner          = 3;
slave_timing[2][64+13].info_temp__j__       = 125;
slave_timing[2][64+13].info_i__quite_rec__  = 0.003000000;
slave_timing[2][64+13].info_dtr__ib__       = -1;
slave_timing[2][64+13].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+13].info_i__max_slave__  = 0.025000000;
slave_timing[2][64+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][64+13].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+13].t_rxd1[0][1] = 2295ns;
slave_timing[2][64+13].t_rxd1[1][0] = 2353ns;
slave_timing[2][64+13].t_rxd1[0][2] = 1749ns;
slave_timing[2][64+13].t_rxd1[2][0] = 2812ns;
slave_timing[2][64+13].t_rxd2[0][2] = 2485ns;
slave_timing[2][64+13].t_rxd2[2][0] = 1787ns;
slave_timing[2][64+13].t_rxd2[1][2] = 1987ns;
slave_timing[2][64+13].t_rxd2[2][1] = 2382ns;

slave_timing[2][64+14].info_corner          = 3;
slave_timing[2][64+14].info_temp__j__       = 125;
slave_timing[2][64+14].info_i__quite_rec__  = 0.003000000;
slave_timing[2][64+14].info_dtr__ib__       = 1;
slave_timing[2][64+14].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+14].info_i__max_slave__  = 0.023000000;
slave_timing[2][64+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][64+14].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+14].t_rxd1[0][1] = 2414ns;
slave_timing[2][64+14].t_rxd1[1][0] = 2196ns;
slave_timing[2][64+14].t_rxd1[0][2] = 1823ns;
slave_timing[2][64+14].t_rxd1[2][0] = 2673ns;
slave_timing[2][64+14].t_rxd2[0][2] = 2764ns;
slave_timing[2][64+14].t_rxd2[2][0] = 1542ns;
slave_timing[2][64+14].t_rxd2[1][2] = 2388ns;
slave_timing[2][64+14].t_rxd2[2][1] = 1960ns;

slave_timing[2][64+15].info_corner          = 3;
slave_timing[2][64+15].info_temp__j__       = 125;
slave_timing[2][64+15].info_i__quite_rec__  = 0.003000000;
slave_timing[2][64+15].info_dtr__ib__       = 1;
slave_timing[2][64+15].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+15].info_i__max_slave__  = 0.025000000;
slave_timing[2][64+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][64+15].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+15].t_rxd1[0][1] = 2310ns;
slave_timing[2][64+15].t_rxd1[1][0] = 2260ns;
slave_timing[2][64+15].t_rxd1[0][2] = 1771ns;
slave_timing[2][64+15].t_rxd1[2][0] = 2714ns;
slave_timing[2][64+15].t_rxd2[0][2] = 2588ns;
slave_timing[2][64+15].t_rxd2[2][0] = 1677ns;
slave_timing[2][64+15].t_rxd2[1][2] = 2142ns;
slave_timing[2][64+15].t_rxd2[2][1] = 2196ns;

slave_timing[2][64+16].info_corner          = 3;
slave_timing[2][64+16].info_temp__j__       = 125;
slave_timing[2][64+16].info_i__quite_rec__  = 0.000000000;
slave_timing[2][64+16].info_dtr__ib__       = -1;
slave_timing[2][64+16].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+16].info_i__max_slave__  = 0.023000000;
slave_timing[2][64+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][64+16].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+16].t_rxd1[0][1] = 2101ns;
slave_timing[2][64+16].t_rxd1[1][0] = 2123ns;
slave_timing[2][64+16].t_rxd1[0][2] = 1604ns;
slave_timing[2][64+16].t_rxd1[2][0] = 2567ns;
slave_timing[2][64+16].t_rxd2[0][2] = 2568ns;
slave_timing[2][64+16].t_rxd2[2][0] = 1611ns;
slave_timing[2][64+16].t_rxd2[1][2] = 2142ns;
slave_timing[2][64+16].t_rxd2[2][1] = 2124ns;

slave_timing[2][64+17].info_corner          = 3;
slave_timing[2][64+17].info_temp__j__       = 125;
slave_timing[2][64+17].info_i__quite_rec__  = 0.000000000;
slave_timing[2][64+17].info_dtr__ib__       = -1;
slave_timing[2][64+17].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+17].info_i__max_slave__  = 0.025000000;
slave_timing[2][64+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][64+17].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+17].t_rxd1[0][1] = 2040ns;
slave_timing[2][64+17].t_rxd1[1][0] = 2184ns;
slave_timing[2][64+17].t_rxd1[0][2] = 1558ns;
slave_timing[2][64+17].t_rxd1[2][0] = 2607ns;
slave_timing[2][64+17].t_rxd2[0][2] = 2419ns;
slave_timing[2][64+17].t_rxd2[2][0] = 1726ns;
slave_timing[2][64+17].t_rxd2[1][2] = 1914ns;
slave_timing[2][64+17].t_rxd2[2][1] = 2345ns;

slave_timing[2][64+18].info_corner          = 3;
slave_timing[2][64+18].info_temp__j__       = 125;
slave_timing[2][64+18].info_i__quite_rec__  = 0.000000000;
slave_timing[2][64+18].info_dtr__ib__       = 1;
slave_timing[2][64+18].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+18].info_i__max_slave__  = 0.023000000;
slave_timing[2][64+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][64+18].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+18].t_rxd1[0][1] = 2188ns;
slave_timing[2][64+18].t_rxd1[1][0] = 2021ns;
slave_timing[2][64+18].t_rxd1[0][2] = 1637ns;
slave_timing[2][64+18].t_rxd1[2][0] = 2498ns;
slave_timing[2][64+18].t_rxd2[0][2] = 2708ns;
slave_timing[2][64+18].t_rxd2[2][0] = 1464ns;
slave_timing[2][64+18].t_rxd2[1][2] = 2347ns;
slave_timing[2][64+18].t_rxd2[2][1] = 1906ns;

slave_timing[2][64+19].info_corner          = 3;
slave_timing[2][64+19].info_temp__j__       = 125;
slave_timing[2][64+19].info_i__quite_rec__  = 0.000000000;
slave_timing[2][64+19].info_dtr__ib__       = 1;
slave_timing[2][64+19].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+19].info_i__max_slave__  = 0.025000000;
slave_timing[2][64+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][64+19].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+19].t_rxd1[0][1] = 2105ns;
slave_timing[2][64+19].t_rxd1[1][0] = 2094ns;
slave_timing[2][64+19].t_rxd1[0][2] = 1588ns;
slave_timing[2][64+19].t_rxd1[2][0] = 2534ns;
slave_timing[2][64+19].t_rxd2[0][2] = 2527ns;
slave_timing[2][64+19].t_rxd2[2][0] = 1614ns;
slave_timing[2][64+19].t_rxd2[1][2] = 2087ns;
slave_timing[2][64+19].t_rxd2[2][1] = 2126ns;

slave_timing[2][64+20].info_corner          = 3;
slave_timing[2][64+20].info_temp__j__       = 125;
slave_timing[2][64+20].info_i__quite_rec__  = 0.000000000;
slave_timing[2][64+20].info_dtr__ib__       = -1;
slave_timing[2][64+20].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+20].info_i__max_slave__  = 0.023000000;
slave_timing[2][64+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][64+20].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+20].t_rxd1[0][1] = 2351ns;
slave_timing[2][64+20].t_rxd1[1][0] = 2268ns;
slave_timing[2][64+20].t_rxd1[0][2] = 1800ns;
slave_timing[2][64+20].t_rxd1[2][0] = 2706ns;
slave_timing[2][64+20].t_rxd2[0][2] = 2598ns;
slave_timing[2][64+20].t_rxd2[2][0] = 1644ns;
slave_timing[2][64+20].t_rxd2[1][2] = 2165ns;
slave_timing[2][64+20].t_rxd2[2][1] = 2142ns;

slave_timing[2][64+21].info_corner          = 3;
slave_timing[2][64+21].info_temp__j__       = 125;
slave_timing[2][64+21].info_i__quite_rec__  = 0.000000000;
slave_timing[2][64+21].info_dtr__ib__       = -1;
slave_timing[2][64+21].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+21].info_i__max_slave__  = 0.025000000;
slave_timing[2][64+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][64+21].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+21].t_rxd1[0][1] = 2270ns;
slave_timing[2][64+21].t_rxd1[1][0] = 2336ns;
slave_timing[2][64+21].t_rxd1[0][2] = 1750ns;
slave_timing[2][64+21].t_rxd1[2][0] = 2746ns;
slave_timing[2][64+21].t_rxd2[0][2] = 2451ns;
slave_timing[2][64+21].t_rxd2[2][0] = 1755ns;
slave_timing[2][64+21].t_rxd2[1][2] = 1941ns;
slave_timing[2][64+21].t_rxd2[2][1] = 2366ns;

slave_timing[2][64+22].info_corner          = 3;
slave_timing[2][64+22].info_temp__j__       = 125;
slave_timing[2][64+22].info_i__quite_rec__  = 0.000000000;
slave_timing[2][64+22].info_dtr__ib__       = 1;
slave_timing[2][64+22].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+22].info_i__max_slave__  = 0.023000000;
slave_timing[2][64+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][64+22].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+22].t_rxd1[0][1] = 2410ns;
slave_timing[2][64+22].t_rxd1[1][0] = 2163ns;
slave_timing[2][64+22].t_rxd1[0][2] = 1826ns;
slave_timing[2][64+22].t_rxd1[2][0] = 2630ns;
slave_timing[2][64+22].t_rxd2[0][2] = 2726ns;
slave_timing[2][64+22].t_rxd2[2][0] = 1511ns;
slave_timing[2][64+22].t_rxd2[1][2] = 2369ns;
slave_timing[2][64+22].t_rxd2[2][1] = 1935ns;

slave_timing[2][64+23].info_corner          = 3;
slave_timing[2][64+23].info_temp__j__       = 125;
slave_timing[2][64+23].info_i__quite_rec__  = 0.000000000;
slave_timing[2][64+23].info_dtr__ib__       = 1;
slave_timing[2][64+23].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+23].info_i__max_slave__  = 0.025000000;
slave_timing[2][64+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][64+23].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+23].t_rxd1[0][1] = 2318ns;
slave_timing[2][64+23].t_rxd1[1][0] = 2235ns;
slave_timing[2][64+23].t_rxd1[0][2] = 1774ns;
slave_timing[2][64+23].t_rxd1[2][0] = 2669ns;
slave_timing[2][64+23].t_rxd2[0][2] = 2545ns;
slave_timing[2][64+23].t_rxd2[2][0] = 1641ns;
slave_timing[2][64+23].t_rxd2[1][2] = 2124ns;
slave_timing[2][64+23].t_rxd2[2][1] = 2154ns;

slave_timing[2][64+24].info_corner          = 3;
slave_timing[2][64+24].info_temp__j__       = 125;
slave_timing[2][64+24].info_i__quite_rec__  = 0.040000000;
slave_timing[2][64+24].info_dtr__ib__       = -1;
slave_timing[2][64+24].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+24].info_i__max_slave__  = 0.023000000;
slave_timing[2][64+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][64+24].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+24].t_rxd1[0][1] = 2204ns;
slave_timing[2][64+24].t_rxd1[1][0] = 2219ns;
slave_timing[2][64+24].t_rxd1[0][2] = 1671ns;
slave_timing[2][64+24].t_rxd1[2][0] = 2688ns;
slave_timing[2][64+24].t_rxd2[0][2] = 2670ns;
slave_timing[2][64+24].t_rxd2[2][0] = 1676ns;
slave_timing[2][64+24].t_rxd2[1][2] = 2197ns;
slave_timing[2][64+24].t_rxd2[2][1] = 2182ns;

slave_timing[2][64+25].info_corner          = 3;
slave_timing[2][64+25].info_temp__j__       = 125;
slave_timing[2][64+25].info_i__quite_rec__  = 0.040000000;
slave_timing[2][64+25].info_dtr__ib__       = -1;
slave_timing[2][64+25].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+25].info_i__max_slave__  = 0.025000000;
slave_timing[2][64+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][64+25].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+25].t_rxd1[0][1] = 2121ns;
slave_timing[2][64+25].t_rxd1[1][0] = 2282ns;
slave_timing[2][64+25].t_rxd1[0][2] = 1627ns;
slave_timing[2][64+25].t_rxd1[2][0] = 2734ns;
slave_timing[2][64+25].t_rxd2[0][2] = 2528ns;
slave_timing[2][64+25].t_rxd2[2][0] = 1801ns;
slave_timing[2][64+25].t_rxd2[1][2] = 1965ns;
slave_timing[2][64+25].t_rxd2[2][1] = 2417ns;

slave_timing[2][64+26].info_corner          = 3;
slave_timing[2][64+26].info_temp__j__       = 125;
slave_timing[2][64+26].info_i__quite_rec__  = 0.040000000;
slave_timing[2][64+26].info_dtr__ib__       = 1;
slave_timing[2][64+26].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+26].info_i__max_slave__  = 0.023000000;
slave_timing[2][64+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][64+26].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+26].t_rxd1[0][1] = 2267ns;
slave_timing[2][64+26].t_rxd1[1][0] = 2164ns;
slave_timing[2][64+26].t_rxd1[0][2] = 1706ns;
slave_timing[2][64+26].t_rxd1[2][0] = 2653ns;
slave_timing[2][64+26].t_rxd2[0][2] = 2804ns;
slave_timing[2][64+26].t_rxd2[2][0] = 1586ns;
slave_timing[2][64+26].t_rxd2[1][2] = 2385ns;
slave_timing[2][64+26].t_rxd2[2][1] = 2015ns;

slave_timing[2][64+27].info_corner          = 3;
slave_timing[2][64+27].info_temp__j__       = 125;
slave_timing[2][64+27].info_i__quite_rec__  = 0.040000000;
slave_timing[2][64+27].info_dtr__ib__       = 1;
slave_timing[2][64+27].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+27].info_i__max_slave__  = 0.025000000;
slave_timing[2][64+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][64+27].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+27].t_rxd1[0][1] = 2174ns;
slave_timing[2][64+27].t_rxd1[1][0] = 2240ns;
slave_timing[2][64+27].t_rxd1[0][2] = 1649ns;
slave_timing[2][64+27].t_rxd1[2][0] = 2700ns;
slave_timing[2][64+27].t_rxd2[0][2] = 2639ns;
slave_timing[2][64+27].t_rxd2[2][0] = 1723ns;
slave_timing[2][64+27].t_rxd2[1][2] = 2135ns;
slave_timing[2][64+27].t_rxd2[2][1] = 2255ns;

slave_timing[2][64+28].info_corner          = 3;
slave_timing[2][64+28].info_temp__j__       = 125;
slave_timing[2][64+28].info_i__quite_rec__  = 0.040000000;
slave_timing[2][64+28].info_dtr__ib__       = -1;
slave_timing[2][64+28].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+28].info_i__max_slave__  = 0.023000000;
slave_timing[2][64+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][64+28].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+28].t_rxd1[0][1] = 2293ns;
slave_timing[2][64+28].t_rxd1[1][0] = 2305ns;
slave_timing[2][64+28].t_rxd1[0][2] = 1762ns;
slave_timing[2][64+28].t_rxd1[2][0] = 2648ns;
slave_timing[2][64+28].t_rxd2[0][2] = 2738ns;
slave_timing[2][64+28].t_rxd2[2][0] = 1991ns;
slave_timing[2][64+28].t_rxd2[1][2] = 2264ns;
slave_timing[2][64+28].t_rxd2[2][1] = 2499ns;

slave_timing[2][64+29].info_corner          = 3;
slave_timing[2][64+29].info_temp__j__       = 125;
slave_timing[2][64+29].info_i__quite_rec__  = 0.040000000;
slave_timing[2][64+29].info_dtr__ib__       = -1;
slave_timing[2][64+29].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+29].info_i__max_slave__  = 0.025000000;
slave_timing[2][64+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][64+29].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+29].t_rxd1[0][1] = 2215ns;
slave_timing[2][64+29].t_rxd1[1][0] = 2375ns;
slave_timing[2][64+29].t_rxd1[0][2] = 1718ns;
slave_timing[2][64+29].t_rxd1[2][0] = 2662ns;
slave_timing[2][64+29].t_rxd2[0][2] = 2608ns;
slave_timing[2][64+29].t_rxd2[2][0] = 2161ns;
slave_timing[2][64+29].t_rxd2[1][2] = 2039ns;
slave_timing[2][64+29].t_rxd2[2][1] = 2803ns;

slave_timing[2][64+30].info_corner          = 3;
slave_timing[2][64+30].info_temp__j__       = 125;
slave_timing[2][64+30].info_i__quite_rec__  = 0.040000000;
slave_timing[2][64+30].info_dtr__ib__       = 1;
slave_timing[2][64+30].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+30].info_i__max_slave__  = 0.023000000;
slave_timing[2][64+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][64+30].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+30].t_rxd1[0][1] = 2356ns;
slave_timing[2][64+30].t_rxd1[1][0] = 2248ns;
slave_timing[2][64+30].t_rxd1[0][2] = 1794ns;
slave_timing[2][64+30].t_rxd1[2][0] = 2654ns;
slave_timing[2][64+30].t_rxd2[0][2] = 2875ns;
slave_timing[2][64+30].t_rxd2[2][0] = 1876ns;
slave_timing[2][64+30].t_rxd2[1][2] = 2453ns;
slave_timing[2][64+30].t_rxd2[2][1] = 2323ns;

slave_timing[2][64+31].info_corner          = 3;
slave_timing[2][64+31].info_temp__j__       = 125;
slave_timing[2][64+31].info_i__quite_rec__  = 0.040000000;
slave_timing[2][64+31].info_dtr__ib__       = 1;
slave_timing[2][64+31].info_i__offset_rec__ = 0.000000000;
slave_timing[2][64+31].info_i__max_slave__  = 0.025000000;
slave_timing[2][64+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][64+31].info_r__dsi_bus__    = 5.000;

slave_timing[2][64+31].t_rxd1[0][1] = 2252ns;
slave_timing[2][64+31].t_rxd1[1][0] = 2312ns;
slave_timing[2][64+31].t_rxd1[0][2] = 1744ns;
slave_timing[2][64+31].t_rxd1[2][0] = 2655ns;
slave_timing[2][64+31].t_rxd2[0][2] = 2720ns;
slave_timing[2][64+31].t_rxd2[2][0] = 2065ns;
slave_timing[2][64+31].t_rxd2[1][2] = 2218ns;
slave_timing[2][64+31].t_rxd2[2][1] = 2635ns;

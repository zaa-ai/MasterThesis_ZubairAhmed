/**
 * Interface: OTP_model_if
 * 
 * interface for setting and reading new OTP data files
 */
interface OTP_model_if;

	string dat_file;
	
endinterface



//-----------------------------------------------------------------------------
// Copyright (c) 2023 Elmos SE
// Author     : Eugene - Easy UVM Generator
//
// Description: This file has been generated automatically by Eugene
//				This file should not be modified manually. 
//-----------------------------------------------------------------------------
`ifndef BUFFER_WRITER_MONITOR_SV
`define BUFFER_WRITER_MONITOR_SV

class buffer_writer_monitor extends uvm_monitor;

	`uvm_component_utils(buffer_writer_monitor)
	
	virtual	buffer_writer_if vif;

  	buffer_writer_config m_config;

  	uvm_analysis_port #(buffer_writer_tr) analysis_port;

  	buffer_writer_tr m_trans;

  	function new(string name, uvm_component parent);
  		super.new(name, parent);
  		analysis_port = new("analysis_port", this);
	endfunction
		
	// Methods run_phase, and do_mon generated by setting monitor_inc in file spi.tpl
	task run_phase(uvm_phase phase);
		`uvm_info(get_type_name(), "run_phase", UVM_HIGH)
		m_trans = buffer_writer_tr::type_id::create("m_trans");
		do_mon();
	endtask
	
	`include "includes/buffer_writer_monitor_inc.sv"
	
	`include "includes/buffer_writer_monitor_inc_inside_class.sv"
	
endclass

// You can insert code here by setting monitor_inc_after_class in file buffer_writer.tpl

`endif

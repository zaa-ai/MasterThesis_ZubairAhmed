
slave_timing[0][96+0].info_corner          = 4;
slave_timing[0][96+0].info_temp__j__       = 125;
slave_timing[0][96+0].info_i__quite_rec__  = 0.006000000;
slave_timing[0][96+0].info_dtr__ib__       = -1;
slave_timing[0][96+0].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+0].info_i__max_slave__  = 0.023000000;
slave_timing[0][96+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][96+0].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+0].t_rxd1[0][1] = 1086ns;
slave_timing[0][96+0].t_rxd1[1][0] = 1089ns;
slave_timing[0][96+0].t_rxd1[0][2] = 807ns;
slave_timing[0][96+0].t_rxd1[2][0] = 1347ns;
slave_timing[0][96+0].t_rxd2[0][2] = 1361ns;
slave_timing[0][96+0].t_rxd2[2][0] = 821ns;
slave_timing[0][96+0].t_rxd2[1][2] = 1116ns;
slave_timing[0][96+0].t_rxd2[2][1] = 1088ns;

slave_timing[0][96+1].info_corner          = 4;
slave_timing[0][96+1].info_temp__j__       = 125;
slave_timing[0][96+1].info_i__quite_rec__  = 0.006000000;
slave_timing[0][96+1].info_dtr__ib__       = -1;
slave_timing[0][96+1].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+1].info_i__max_slave__  = 0.025000000;
slave_timing[0][96+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][96+1].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+1].t_rxd1[0][1] = 1040ns;
slave_timing[0][96+1].t_rxd1[1][0] = 1117ns;
slave_timing[0][96+1].t_rxd1[0][2] = 784ns;
slave_timing[0][96+1].t_rxd1[2][0] = 1375ns;
slave_timing[0][96+1].t_rxd2[0][2] = 1259ns;
slave_timing[0][96+1].t_rxd2[2][0] = 874ns;
slave_timing[0][96+1].t_rxd2[1][2] = 991ns;
slave_timing[0][96+1].t_rxd2[2][1] = 1212ns;

slave_timing[0][96+2].info_corner          = 4;
slave_timing[0][96+2].info_temp__j__       = 125;
slave_timing[0][96+2].info_i__quite_rec__  = 0.006000000;
slave_timing[0][96+2].info_dtr__ib__       = 1;
slave_timing[0][96+2].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+2].info_i__max_slave__  = 0.023000000;
slave_timing[0][96+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][96+2].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+2].t_rxd1[0][1] = 1086ns;
slave_timing[0][96+2].t_rxd1[1][0] = 1047ns;
slave_timing[0][96+2].t_rxd1[0][2] = 802ns;
slave_timing[0][96+2].t_rxd1[2][0] = 1297ns;
slave_timing[0][96+2].t_rxd2[0][2] = 1412ns;
slave_timing[0][96+2].t_rxd2[2][0] = 775ns;
slave_timing[0][96+2].t_rxd2[1][2] = 1190ns;
slave_timing[0][96+2].t_rxd2[2][1] = 1003ns;

slave_timing[0][96+3].info_corner          = 4;
slave_timing[0][96+3].info_temp__j__       = 125;
slave_timing[0][96+3].info_i__quite_rec__  = 0.006000000;
slave_timing[0][96+3].info_dtr__ib__       = 1;
slave_timing[0][96+3].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+3].info_i__max_slave__  = 0.025000000;
slave_timing[0][96+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][96+3].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+3].t_rxd1[0][1] = 1039ns;
slave_timing[0][96+3].t_rxd1[1][0] = 1081ns;
slave_timing[0][96+3].t_rxd1[0][2] = 778ns;
slave_timing[0][96+3].t_rxd1[2][0] = 1325ns;
slave_timing[0][96+3].t_rxd2[0][2] = 1290ns;
slave_timing[0][96+3].t_rxd2[2][0] = 831ns;
slave_timing[0][96+3].t_rxd2[1][2] = 1051ns;
slave_timing[0][96+3].t_rxd2[2][1] = 1118ns;

slave_timing[0][96+4].info_corner          = 4;
slave_timing[0][96+4].info_temp__j__       = 125;
slave_timing[0][96+4].info_i__quite_rec__  = 0.006000000;
slave_timing[0][96+4].info_dtr__ib__       = -1;
slave_timing[0][96+4].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+4].info_i__max_slave__  = 0.023000000;
slave_timing[0][96+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][96+4].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+4].t_rxd1[0][1] = 1273ns;
slave_timing[0][96+4].t_rxd1[1][0] = 1220ns;
slave_timing[0][96+4].t_rxd1[0][2] = 934ns;
slave_timing[0][96+4].t_rxd1[2][0] = 1468ns;
slave_timing[0][96+4].t_rxd2[0][2] = 1423ns;
slave_timing[0][96+4].t_rxd2[2][0] = 860ns;
slave_timing[0][96+4].t_rxd2[1][2] = 1140ns;
slave_timing[0][96+4].t_rxd2[2][1] = 1112ns;

slave_timing[0][96+5].info_corner          = 4;
slave_timing[0][96+5].info_temp__j__       = 125;
slave_timing[0][96+5].info_i__quite_rec__  = 0.006000000;
slave_timing[0][96+5].info_dtr__ib__       = -1;
slave_timing[0][96+5].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+5].info_i__max_slave__  = 0.025000000;
slave_timing[0][96+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][96+5].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+5].t_rxd1[0][1] = 1215ns;
slave_timing[0][96+5].t_rxd1[1][0] = 1251ns;
slave_timing[0][96+5].t_rxd1[0][2] = 907ns;
slave_timing[0][96+5].t_rxd1[2][0] = 1493ns;
slave_timing[0][96+5].t_rxd2[0][2] = 1322ns;
slave_timing[0][96+5].t_rxd2[2][0] = 911ns;
slave_timing[0][96+5].t_rxd2[1][2] = 1018ns;
slave_timing[0][96+5].t_rxd2[2][1] = 1215ns;

slave_timing[0][96+6].info_corner          = 4;
slave_timing[0][96+6].info_temp__j__       = 125;
slave_timing[0][96+6].info_i__quite_rec__  = 0.006000000;
slave_timing[0][96+6].info_dtr__ib__       = 1;
slave_timing[0][96+6].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+6].info_i__max_slave__  = 0.023000000;
slave_timing[0][96+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][96+6].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+6].t_rxd1[0][1] = 1273ns;
slave_timing[0][96+6].t_rxd1[1][0] = 1171ns;
slave_timing[0][96+6].t_rxd1[0][2] = 928ns;
slave_timing[0][96+6].t_rxd1[2][0] = 1411ns;
slave_timing[0][96+6].t_rxd2[0][2] = 1468ns;
slave_timing[0][96+6].t_rxd2[2][0] = 809ns;
slave_timing[0][96+6].t_rxd2[1][2] = 1210ns;
slave_timing[0][96+6].t_rxd2[2][1] = 1025ns;

slave_timing[0][96+7].info_corner          = 4;
slave_timing[0][96+7].info_temp__j__       = 125;
slave_timing[0][96+7].info_i__quite_rec__  = 0.006000000;
slave_timing[0][96+7].info_dtr__ib__       = 1;
slave_timing[0][96+7].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+7].info_i__max_slave__  = 0.025000000;
slave_timing[0][96+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][96+7].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+7].t_rxd1[0][1] = 1213ns;
slave_timing[0][96+7].t_rxd1[1][0] = 1201ns;
slave_timing[0][96+7].t_rxd1[0][2] = 901ns;
slave_timing[0][96+7].t_rxd1[2][0] = 1436ns;
slave_timing[0][96+7].t_rxd2[0][2] = 1349ns;
slave_timing[0][96+7].t_rxd2[2][0] = 865ns;
slave_timing[0][96+7].t_rxd2[1][2] = 1074ns;
slave_timing[0][96+7].t_rxd2[2][1] = 1126ns;

slave_timing[0][96+8].info_corner          = 4;
slave_timing[0][96+8].info_temp__j__       = 125;
slave_timing[0][96+8].info_i__quite_rec__  = 0.003000000;
slave_timing[0][96+8].info_dtr__ib__       = -1;
slave_timing[0][96+8].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+8].info_i__max_slave__  = 0.023000000;
slave_timing[0][96+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][96+8].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+8].t_rxd1[0][1] = 1052ns;
slave_timing[0][96+8].t_rxd1[1][0] = 1056ns;
slave_timing[0][96+8].t_rxd1[0][2] = 785ns;
slave_timing[0][96+8].t_rxd1[2][0] = 1293ns;
slave_timing[0][96+8].t_rxd2[0][2] = 1309ns;
slave_timing[0][96+8].t_rxd2[2][0] = 802ns;
slave_timing[0][96+8].t_rxd2[1][2] = 1089ns;
slave_timing[0][96+8].t_rxd2[2][1] = 1055ns;

slave_timing[0][96+9].info_corner          = 4;
slave_timing[0][96+9].info_temp__j__       = 125;
slave_timing[0][96+9].info_i__quite_rec__  = 0.003000000;
slave_timing[0][96+9].info_dtr__ib__       = -1;
slave_timing[0][96+9].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+9].info_i__max_slave__  = 0.025000000;
slave_timing[0][96+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][96+9].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+9].t_rxd1[0][1] = 1006ns;
slave_timing[0][96+9].t_rxd1[1][0] = 1083ns;
slave_timing[0][96+9].t_rxd1[0][2] = 762ns;
slave_timing[0][96+9].t_rxd1[2][0] = 1317ns;
slave_timing[0][96+9].t_rxd2[0][2] = 1213ns;
slave_timing[0][96+9].t_rxd2[2][0] = 854ns;
slave_timing[0][96+9].t_rxd2[1][2] = 968ns;
slave_timing[0][96+9].t_rxd2[2][1] = 1173ns;

slave_timing[0][96+10].info_corner          = 4;
slave_timing[0][96+10].info_temp__j__       = 125;
slave_timing[0][96+10].info_i__quite_rec__  = 0.003000000;
slave_timing[0][96+10].info_dtr__ib__       = 1;
slave_timing[0][96+10].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+10].info_i__max_slave__  = 0.023000000;
slave_timing[0][96+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][96+10].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+10].t_rxd1[0][1] = 1060ns;
slave_timing[0][96+10].t_rxd1[1][0] = 1022ns;
slave_timing[0][96+10].t_rxd1[0][2] = 785ns;
slave_timing[0][96+10].t_rxd1[2][0] = 1245ns;
slave_timing[0][96+10].t_rxd2[0][2] = 1356ns;
slave_timing[0][96+10].t_rxd2[2][0] = 746ns;
slave_timing[0][96+10].t_rxd2[1][2] = 1158ns;
slave_timing[0][96+10].t_rxd2[2][1] = 962ns;

slave_timing[0][96+11].info_corner          = 4;
slave_timing[0][96+11].info_temp__j__       = 125;
slave_timing[0][96+11].info_i__quite_rec__  = 0.003000000;
slave_timing[0][96+11].info_dtr__ib__       = 1;
slave_timing[0][96+11].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+11].info_i__max_slave__  = 0.025000000;
slave_timing[0][96+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][96+11].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+11].t_rxd1[0][1] = 1013ns;
slave_timing[0][96+11].t_rxd1[1][0] = 1051ns;
slave_timing[0][96+11].t_rxd1[0][2] = 760ns;
slave_timing[0][96+11].t_rxd1[2][0] = 1268ns;
slave_timing[0][96+11].t_rxd2[0][2] = 1240ns;
slave_timing[0][96+11].t_rxd2[2][0] = 803ns;
slave_timing[0][96+11].t_rxd2[1][2] = 1021ns;
slave_timing[0][96+11].t_rxd2[2][1] = 1070ns;

slave_timing[0][96+12].info_corner          = 4;
slave_timing[0][96+12].info_temp__j__       = 125;
slave_timing[0][96+12].info_i__quite_rec__  = 0.003000000;
slave_timing[0][96+12].info_dtr__ib__       = -1;
slave_timing[0][96+12].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+12].info_i__max_slave__  = 0.023000000;
slave_timing[0][96+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][96+12].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+12].t_rxd1[0][1] = 1254ns;
slave_timing[0][96+12].t_rxd1[1][0] = 1185ns;
slave_timing[0][96+12].t_rxd1[0][2] = 923ns;
slave_timing[0][96+12].t_rxd1[2][0] = 1409ns;
slave_timing[0][96+12].t_rxd2[0][2] = 1371ns;
slave_timing[0][96+12].t_rxd2[2][0] = 837ns;
slave_timing[0][96+12].t_rxd2[1][2] = 1107ns;
slave_timing[0][96+12].t_rxd2[2][1] = 1069ns;

slave_timing[0][96+13].info_corner          = 4;
slave_timing[0][96+13].info_temp__j__       = 125;
slave_timing[0][96+13].info_i__quite_rec__  = 0.003000000;
slave_timing[0][96+13].info_dtr__ib__       = -1;
slave_timing[0][96+13].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+13].info_i__max_slave__  = 0.025000000;
slave_timing[0][96+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][96+13].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+13].t_rxd1[0][1] = 1198ns;
slave_timing[0][96+13].t_rxd1[1][0] = 1213ns;
slave_timing[0][96+13].t_rxd1[0][2] = 897ns;
slave_timing[0][96+13].t_rxd1[2][0] = 1433ns;
slave_timing[0][96+13].t_rxd2[0][2] = 1278ns;
slave_timing[0][96+13].t_rxd2[2][0] = 888ns;
slave_timing[0][96+13].t_rxd2[1][2] = 995ns;
slave_timing[0][96+13].t_rxd2[2][1] = 1189ns;

slave_timing[0][96+14].info_corner          = 4;
slave_timing[0][96+14].info_temp__j__       = 125;
slave_timing[0][96+14].info_i__quite_rec__  = 0.003000000;
slave_timing[0][96+14].info_dtr__ib__       = 1;
slave_timing[0][96+14].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+14].info_i__max_slave__  = 0.023000000;
slave_timing[0][96+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][96+14].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+14].t_rxd1[0][1] = 1262ns;
slave_timing[0][96+14].t_rxd1[1][0] = 1143ns;
slave_timing[0][96+14].t_rxd1[0][2] = 922ns;
slave_timing[0][96+14].t_rxd1[2][0] = 1357ns;
slave_timing[0][96+14].t_rxd2[0][2] = 1413ns;
slave_timing[0][96+14].t_rxd2[2][0] = 781ns;
slave_timing[0][96+14].t_rxd2[1][2] = 1175ns;
slave_timing[0][96+14].t_rxd2[2][1] = 987ns;

slave_timing[0][96+15].info_corner          = 4;
slave_timing[0][96+15].info_temp__j__       = 125;
slave_timing[0][96+15].info_i__quite_rec__  = 0.003000000;
slave_timing[0][96+15].info_dtr__ib__       = 1;
slave_timing[0][96+15].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+15].info_i__max_slave__  = 0.025000000;
slave_timing[0][96+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][96+15].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+15].t_rxd1[0][1] = 1203ns;
slave_timing[0][96+15].t_rxd1[1][0] = 1173ns;
slave_timing[0][96+15].t_rxd1[0][2] = 894ns;
slave_timing[0][96+15].t_rxd1[2][0] = 1379ns;
slave_timing[0][96+15].t_rxd2[0][2] = 1300ns;
slave_timing[0][96+15].t_rxd2[2][0] = 837ns;
slave_timing[0][96+15].t_rxd2[1][2] = 1043ns;
slave_timing[0][96+15].t_rxd2[2][1] = 1090ns;

slave_timing[0][96+16].info_corner          = 4;
slave_timing[0][96+16].info_temp__j__       = 125;
slave_timing[0][96+16].info_i__quite_rec__  = 0.000000000;
slave_timing[0][96+16].info_dtr__ib__       = -1;
slave_timing[0][96+16].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+16].info_i__max_slave__  = 0.023000000;
slave_timing[0][96+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][96+16].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+16].t_rxd1[0][1] = 1030ns;
slave_timing[0][96+16].t_rxd1[1][0] = 1025ns;
slave_timing[0][96+16].t_rxd1[0][2] = 770ns;
slave_timing[0][96+16].t_rxd1[2][0] = 1235ns;
slave_timing[0][96+16].t_rxd2[0][2] = 1255ns;
slave_timing[0][96+16].t_rxd2[2][0] = 772ns;
slave_timing[0][96+16].t_rxd2[1][2] = 1052ns;
slave_timing[0][96+16].t_rxd2[2][1] = 1013ns;

slave_timing[0][96+17].info_corner          = 4;
slave_timing[0][96+17].info_temp__j__       = 125;
slave_timing[0][96+17].info_i__quite_rec__  = 0.000000000;
slave_timing[0][96+17].info_dtr__ib__       = -1;
slave_timing[0][96+17].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+17].info_i__max_slave__  = 0.025000000;
slave_timing[0][96+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][96+17].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+17].t_rxd1[0][1] = 989ns;
slave_timing[0][96+17].t_rxd1[1][0] = 1052ns;
slave_timing[0][96+17].t_rxd1[0][2] = 747ns;
slave_timing[0][96+17].t_rxd1[2][0] = 1259ns;
slave_timing[0][96+17].t_rxd2[0][2] = 1165ns;
slave_timing[0][96+17].t_rxd2[2][0] = 822ns;
slave_timing[0][96+17].t_rxd2[1][2] = 939ns;
slave_timing[0][96+17].t_rxd2[2][1] = 1122ns;

slave_timing[0][96+18].info_corner          = 4;
slave_timing[0][96+18].info_temp__j__       = 125;
slave_timing[0][96+18].info_i__quite_rec__  = 0.000000000;
slave_timing[0][96+18].info_dtr__ib__       = 1;
slave_timing[0][96+18].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+18].info_i__max_slave__  = 0.023000000;
slave_timing[0][96+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][96+18].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+18].t_rxd1[0][1] = 1036ns;
slave_timing[0][96+18].t_rxd1[1][0] = 987ns;
slave_timing[0][96+18].t_rxd1[0][2] = 767ns;
slave_timing[0][96+18].t_rxd1[2][0] = 1198ns;
slave_timing[0][96+18].t_rxd2[0][2] = 1302ns;
slave_timing[0][96+18].t_rxd2[2][0] = 724ns;
slave_timing[0][96+18].t_rxd2[1][2] = 1116ns;
slave_timing[0][96+18].t_rxd2[2][1] = 926ns;

slave_timing[0][96+19].info_corner          = 4;
slave_timing[0][96+19].info_temp__j__       = 125;
slave_timing[0][96+19].info_i__quite_rec__  = 0.000000000;
slave_timing[0][96+19].info_dtr__ib__       = 1;
slave_timing[0][96+19].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+19].info_i__max_slave__  = 0.025000000;
slave_timing[0][96+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][96+19].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+19].t_rxd1[0][1] = 992ns;
slave_timing[0][96+19].t_rxd1[1][0] = 1018ns;
slave_timing[0][96+19].t_rxd1[0][2] = 745ns;
slave_timing[0][96+19].t_rxd1[2][0] = 1222ns;
slave_timing[0][96+19].t_rxd2[0][2] = 1195ns;
slave_timing[0][96+19].t_rxd2[2][0] = 779ns;
slave_timing[0][96+19].t_rxd2[1][2] = 990ns;
slave_timing[0][96+19].t_rxd2[2][1] = 1031ns;

slave_timing[0][96+20].info_corner          = 4;
slave_timing[0][96+20].info_temp__j__       = 125;
slave_timing[0][96+20].info_i__quite_rec__  = 0.000000000;
slave_timing[0][96+20].info_dtr__ib__       = -1;
slave_timing[0][96+20].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+20].info_i__max_slave__  = 0.023000000;
slave_timing[0][96+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][96+20].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+20].t_rxd1[0][1] = 1257ns;
slave_timing[0][96+20].t_rxd1[1][0] = 1150ns;
slave_timing[0][96+20].t_rxd1[0][2] = 924ns;
slave_timing[0][96+20].t_rxd1[2][0] = 1343ns;
slave_timing[0][96+20].t_rxd2[0][2] = 1315ns;
slave_timing[0][96+20].t_rxd2[2][0] = 807ns;
slave_timing[0][96+20].t_rxd2[1][2] = 1071ns;
slave_timing[0][96+20].t_rxd2[2][1] = 1024ns;

slave_timing[0][96+21].info_corner          = 4;
slave_timing[0][96+21].info_temp__j__       = 125;
slave_timing[0][96+21].info_i__quite_rec__  = 0.000000000;
slave_timing[0][96+21].info_dtr__ib__       = -1;
slave_timing[0][96+21].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+21].info_i__max_slave__  = 0.025000000;
slave_timing[0][96+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][96+21].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+21].t_rxd1[0][1] = 1202ns;
slave_timing[0][96+21].t_rxd1[1][0] = 1175ns;
slave_timing[0][96+21].t_rxd1[0][2] = 896ns;
slave_timing[0][96+21].t_rxd1[2][0] = 1366ns;
slave_timing[0][96+21].t_rxd2[0][2] = 1228ns;
slave_timing[0][96+21].t_rxd2[2][0] = 856ns;
slave_timing[0][96+21].t_rxd2[1][2] = 964ns;
slave_timing[0][96+21].t_rxd2[2][1] = 1137ns;

slave_timing[0][96+22].info_corner          = 4;
slave_timing[0][96+22].info_temp__j__       = 125;
slave_timing[0][96+22].info_i__quite_rec__  = 0.000000000;
slave_timing[0][96+22].info_dtr__ib__       = 1;
slave_timing[0][96+22].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+22].info_i__max_slave__  = 0.023000000;
slave_timing[0][96+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][96+22].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+22].t_rxd1[0][1] = 1262ns;
slave_timing[0][96+22].t_rxd1[1][0] = 1108ns;
slave_timing[0][96+22].t_rxd1[0][2] = 920ns;
slave_timing[0][96+22].t_rxd1[2][0] = 1306ns;
slave_timing[0][96+22].t_rxd2[0][2] = 1357ns;
slave_timing[0][96+22].t_rxd2[2][0] = 758ns;
slave_timing[0][96+22].t_rxd2[1][2] = 1131ns;
slave_timing[0][96+22].t_rxd2[2][1] = 942ns;

slave_timing[0][96+23].info_corner          = 4;
slave_timing[0][96+23].info_temp__j__       = 125;
slave_timing[0][96+23].info_i__quite_rec__  = 0.000000000;
slave_timing[0][96+23].info_dtr__ib__       = 1;
slave_timing[0][96+23].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+23].info_i__max_slave__  = 0.025000000;
slave_timing[0][96+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][96+23].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+23].t_rxd1[0][1] = 1203ns;
slave_timing[0][96+23].t_rxd1[1][0] = 1139ns;
slave_timing[0][96+23].t_rxd1[0][2] = 894ns;
slave_timing[0][96+23].t_rxd1[2][0] = 1328ns;
slave_timing[0][96+23].t_rxd2[0][2] = 1254ns;
slave_timing[0][96+23].t_rxd2[2][0] = 810ns;
slave_timing[0][96+23].t_rxd2[1][2] = 1012ns;
slave_timing[0][96+23].t_rxd2[2][1] = 1039ns;

slave_timing[0][96+24].info_corner          = 4;
slave_timing[0][96+24].info_temp__j__       = 125;
slave_timing[0][96+24].info_i__quite_rec__  = 0.040000000;
slave_timing[0][96+24].info_dtr__ib__       = -1;
slave_timing[0][96+24].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+24].info_i__max_slave__  = 0.023000000;
slave_timing[0][96+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][96+24].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+24].t_rxd1[0][1] = 1175ns;
slave_timing[0][96+24].t_rxd1[1][0] = 1163ns;
slave_timing[0][96+24].t_rxd1[0][2] = 904ns;
slave_timing[0][96+24].t_rxd1[2][0] = 1517ns;
slave_timing[0][96+24].t_rxd2[0][2] = 1660ns;
slave_timing[0][96+24].t_rxd2[2][0] = 1001ns;
slave_timing[0][96+24].t_rxd2[1][2] = 1386ns;
slave_timing[0][96+24].t_rxd2[2][1] = 1344ns;

slave_timing[0][96+25].info_corner          = 4;
slave_timing[0][96+25].info_temp__j__       = 125;
slave_timing[0][96+25].info_i__quite_rec__  = 0.040000000;
slave_timing[0][96+25].info_dtr__ib__       = -1;
slave_timing[0][96+25].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+25].info_i__max_slave__  = 0.025000000;
slave_timing[0][96+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][96+25].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+25].t_rxd1[0][1] = 1132ns;
slave_timing[0][96+25].t_rxd1[1][0] = 1207ns;
slave_timing[0][96+25].t_rxd1[0][2] = 881ns;
slave_timing[0][96+25].t_rxd1[2][0] = 1556ns;
slave_timing[0][96+25].t_rxd2[0][2] = 1541ns;
slave_timing[0][96+25].t_rxd2[2][0] = 1061ns;
slave_timing[0][96+25].t_rxd2[1][2] = 1235ns;
slave_timing[0][96+25].t_rxd2[2][1] = 1503ns;

slave_timing[0][96+26].info_corner          = 4;
slave_timing[0][96+26].info_temp__j__       = 125;
slave_timing[0][96+26].info_i__quite_rec__  = 0.040000000;
slave_timing[0][96+26].info_dtr__ib__       = 1;
slave_timing[0][96+26].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+26].info_i__max_slave__  = 0.023000000;
slave_timing[0][96+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][96+26].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+26].t_rxd1[0][1] = 1209ns;
slave_timing[0][96+26].t_rxd1[1][0] = 1127ns;
slave_timing[0][96+26].t_rxd1[0][2] = 918ns;
slave_timing[0][96+26].t_rxd1[2][0] = 1484ns;
slave_timing[0][96+26].t_rxd2[0][2] = 1763ns;
slave_timing[0][96+26].t_rxd2[2][0] = 949ns;
slave_timing[0][96+26].t_rxd2[1][2] = 1511ns;
slave_timing[0][96+26].t_rxd2[2][1] = 1235ns;

slave_timing[0][96+27].info_corner          = 4;
slave_timing[0][96+27].info_temp__j__       = 125;
slave_timing[0][96+27].info_i__quite_rec__  = 0.040000000;
slave_timing[0][96+27].info_dtr__ib__       = 1;
slave_timing[0][96+27].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+27].info_i__max_slave__  = 0.025000000;
slave_timing[0][96+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][96+27].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+27].t_rxd1[0][1] = 1160ns;
slave_timing[0][96+27].t_rxd1[1][0] = 1171ns;
slave_timing[0][96+27].t_rxd1[0][2] = 893ns;
slave_timing[0][96+27].t_rxd1[2][0] = 1523ns;
slave_timing[0][96+27].t_rxd2[0][2] = 1614ns;
slave_timing[0][96+27].t_rxd2[2][0] = 1014ns;
slave_timing[0][96+27].t_rxd2[1][2] = 1333ns;
slave_timing[0][96+27].t_rxd2[2][1] = 1383ns;

slave_timing[0][96+28].info_corner          = 4;
slave_timing[0][96+28].info_temp__j__       = 125;
slave_timing[0][96+28].info_i__quite_rec__  = 0.040000000;
slave_timing[0][96+28].info_dtr__ib__       = -1;
slave_timing[0][96+28].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+28].info_i__max_slave__  = 0.023000000;
slave_timing[0][96+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][96+28].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+28].t_rxd1[0][1] = 1290ns;
slave_timing[0][96+28].t_rxd1[1][0] = 1603ns;
slave_timing[0][96+28].t_rxd1[0][2] = 1034ns;
slave_timing[0][96+28].t_rxd1[2][0] = 2448ns;
slave_timing[0][96+28].t_rxd2[0][2] = 2590ns;
slave_timing[0][96+28].t_rxd2[2][0] = 1479ns;
slave_timing[0][96+28].t_rxd2[1][2] = 2211ns;
slave_timing[0][96+28].t_rxd2[2][1] = 2193ns;

slave_timing[0][96+29].info_corner          = 4;
slave_timing[0][96+29].info_temp__j__       = 125;
slave_timing[0][96+29].info_i__quite_rec__  = 0.040000000;
slave_timing[0][96+29].info_dtr__ib__       = -1;
slave_timing[0][96+29].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+29].info_i__max_slave__  = 0.025000000;
slave_timing[0][96+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][96+29].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+29].t_rxd1[0][1] = 1251ns;
slave_timing[0][96+29].t_rxd1[1][0] = 1694ns;
slave_timing[0][96+29].t_rxd1[0][2] = 1011ns;
slave_timing[0][96+29].t_rxd1[2][0] = 2554ns;
slave_timing[0][96+29].t_rxd2[0][2] = 2329ns;
slave_timing[0][96+29].t_rxd2[2][0] = 1609ns;
slave_timing[0][96+29].t_rxd2[1][2] = 1883ns;
slave_timing[0][96+29].t_rxd2[2][1] = 2587ns;

slave_timing[0][96+30].info_corner          = 4;
slave_timing[0][96+30].info_temp__j__       = 125;
slave_timing[0][96+30].info_i__quite_rec__  = 0.040000000;
slave_timing[0][96+30].info_dtr__ib__       = 1;
slave_timing[0][96+30].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+30].info_i__max_slave__  = 0.023000000;
slave_timing[0][96+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][96+30].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+30].t_rxd1[0][1] = 1318ns;
slave_timing[0][96+30].t_rxd1[1][0] = 1497ns;
slave_timing[0][96+30].t_rxd1[0][2] = 1030ns;
slave_timing[0][96+30].t_rxd1[2][0] = 2326ns;
slave_timing[0][96+30].t_rxd2[0][2] = 2818ns;
slave_timing[0][96+30].t_rxd2[2][0] = 1379ns;
slave_timing[0][96+30].t_rxd2[1][2] = 2491ns;
slave_timing[0][96+30].t_rxd2[2][1] = 1933ns;

slave_timing[0][96+31].info_corner          = 4;
slave_timing[0][96+31].info_temp__j__       = 125;
slave_timing[0][96+31].info_i__quite_rec__  = 0.040000000;
slave_timing[0][96+31].info_dtr__ib__       = 1;
slave_timing[0][96+31].info_i__offset_rec__ = 0.000000000;
slave_timing[0][96+31].info_i__max_slave__  = 0.025000000;
slave_timing[0][96+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][96+31].info_r__dsi_bus__    = 5.000;

slave_timing[0][96+31].t_rxd1[0][1] = 1272ns;
slave_timing[0][96+31].t_rxd1[1][0] = 1588ns;
slave_timing[0][96+31].t_rxd1[0][2] = 1021ns;
slave_timing[0][96+31].t_rxd1[2][0] = 2427ns;
slave_timing[0][96+31].t_rxd2[0][2] = 2480ns;
slave_timing[0][96+31].t_rxd2[2][0] = 1508ns;
slave_timing[0][96+31].t_rxd2[1][2] = 2088ns;
slave_timing[0][96+31].t_rxd2[2][1] = 2279ns;

/* ###   interface instances   ###################################################### */

ELIP_test_register_IR_ELIP_RDF_if ELIP_test_register_IR_ELIP_RDF (); 
ELIP_test_register_IR_ELIP_RD_if ELIP_test_register_IR_ELIP_RD (); 
ELIP_test_register_IR_ELIP_RDI_if ELIP_test_register_IR_ELIP_RDI (); 
ELIP_test_register_IR_ELIP_WRF_if ELIP_test_register_IR_ELIP_WRF (); 
ELIP_test_register_IR_ELIP_WR_if ELIP_test_register_IR_ELIP_WR (); 
ELIP_test_register_IR_ELIP_WRI_if ELIP_test_register_IR_ELIP_WRI (); 



slave_timing[1][0].info_corner          = 0;
slave_timing[1][0].info_temp__j__       = 25;
slave_timing[1][0].info_i__quite_rec__  = 0.006000000;
slave_timing[1][0].info_dtr__ib__       = -1;
slave_timing[1][0].info_i__offset_rec__ = -0.001000000;
slave_timing[1][0].info_i__max_slave__  = 0.021000000;
slave_timing[1][0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][0].info_r__dsi_bus__    = 5.000;

slave_timing[1][0].t_rxd1[0][1] = 2167ns;
slave_timing[1][0].t_rxd1[1][0] = 1552ns;
slave_timing[1][0].t_rxd1[0][2] = 1483ns;
slave_timing[1][0].t_rxd1[2][0] = 1962ns;
slave_timing[1][0].t_rxd2[0][2] = 2450ns;
slave_timing[1][0].t_rxd2[2][0] = 1216ns;
slave_timing[1][0].t_rxd2[1][2] = 2189ns;
slave_timing[1][0].t_rxd2[2][1] = 1556ns;

slave_timing[1][1].info_corner          = 0;
slave_timing[1][1].info_temp__j__       = 25;
slave_timing[1][1].info_i__quite_rec__  = 0.006000000;
slave_timing[1][1].info_dtr__ib__       = -1;
slave_timing[1][1].info_i__offset_rec__ = 0.001000000;
slave_timing[1][1].info_i__max_slave__  = 0.021000000;
slave_timing[1][1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][1].info_r__dsi_bus__    = 5.000;

slave_timing[1][1].t_rxd1[0][1] = 1810ns;
slave_timing[1][1].t_rxd1[1][0] = 1822ns;
slave_timing[1][1].t_rxd1[0][2] = 1347ns;
slave_timing[1][1].t_rxd1[2][0] = 2158ns;
slave_timing[1][1].t_rxd2[0][2] = 2152ns;
slave_timing[1][1].t_rxd2[2][0] = 1363ns;
slave_timing[1][1].t_rxd2[1][2] = 1827ns;
slave_timing[1][1].t_rxd2[2][1] = 1829ns;

slave_timing[1][2].info_corner          = 0;
slave_timing[1][2].info_temp__j__       = 25;
slave_timing[1][2].info_i__quite_rec__  = 0.006000000;
slave_timing[1][2].info_dtr__ib__       = -1;
slave_timing[1][2].info_i__offset_rec__ = -0.001000000;
slave_timing[1][2].info_i__max_slave__  = 0.027000000;
slave_timing[1][2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][2].info_r__dsi_bus__    = 5.000;

slave_timing[1][2].t_rxd1[0][1] = 1824ns;
slave_timing[1][2].t_rxd1[1][0] = 1714ns;
slave_timing[1][2].t_rxd1[0][2] = 1351ns;
slave_timing[1][2].t_rxd1[2][0] = 2074ns;
slave_timing[1][2].t_rxd2[0][2] = 1933ns;
slave_timing[1][2].t_rxd2[2][0] = 1466ns;
slave_timing[1][2].t_rxd2[1][2] = 1514ns;
slave_timing[1][2].t_rxd2[2][1] = 2097ns;

slave_timing[1][3].info_corner          = 0;
slave_timing[1][3].info_temp__j__       = 25;
slave_timing[1][3].info_i__quite_rec__  = 0.006000000;
slave_timing[1][3].info_dtr__ib__       = -1;
slave_timing[1][3].info_i__offset_rec__ = 0.001000000;
slave_timing[1][3].info_i__max_slave__  = 0.027000000;
slave_timing[1][3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][3].info_r__dsi_bus__    = 5.000;

slave_timing[1][3].t_rxd1[0][1] = 1627ns;
slave_timing[1][3].t_rxd1[1][0] = 1924ns;
slave_timing[1][3].t_rxd1[0][2] = 1236ns;
slave_timing[1][3].t_rxd1[2][0] = 2237ns;
slave_timing[1][3].t_rxd2[0][2] = 1809ns;
slave_timing[1][3].t_rxd2[2][0] = 1562ns;
slave_timing[1][3].t_rxd2[1][2] = 1323ns;
slave_timing[1][3].t_rxd2[2][1] = 2540ns;

slave_timing[1][4].info_corner          = 0;
slave_timing[1][4].info_temp__j__       = 25;
slave_timing[1][4].info_i__quite_rec__  = 0.006000000;
slave_timing[1][4].info_dtr__ib__       = 1;
slave_timing[1][4].info_i__offset_rec__ = -0.001000000;
slave_timing[1][4].info_i__max_slave__  = 0.021000000;
slave_timing[1][4].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][4].info_r__dsi_bus__    = 5.000;

slave_timing[1][4].t_rxd1[0][1] = 2288ns;
slave_timing[1][4].t_rxd1[1][0] = 1511ns;
slave_timing[1][4].t_rxd1[0][2] = 1514ns;
slave_timing[1][4].t_rxd1[2][0] = 1938ns;
slave_timing[1][4].t_rxd2[0][2] = 2797ns;
slave_timing[1][4].t_rxd2[2][0] = 1133ns;
slave_timing[1][4].t_rxd2[1][2] = 2562ns;
slave_timing[1][4].t_rxd2[2][1] = 1424ns;

slave_timing[1][5].info_corner          = 0;
slave_timing[1][5].info_temp__j__       = 25;
slave_timing[1][5].info_i__quite_rec__  = 0.006000000;
slave_timing[1][5].info_dtr__ib__       = 1;
slave_timing[1][5].info_i__offset_rec__ = 0.001000000;
slave_timing[1][5].info_i__max_slave__  = 0.021000000;
slave_timing[1][5].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][5].info_r__dsi_bus__    = 5.000;

slave_timing[1][5].t_rxd1[0][1] = 1884ns;
slave_timing[1][5].t_rxd1[1][0] = 1780ns;
slave_timing[1][5].t_rxd1[0][2] = 1380ns;
slave_timing[1][5].t_rxd1[2][0] = 2124ns;
slave_timing[1][5].t_rxd2[0][2] = 2303ns;
slave_timing[1][5].t_rxd2[2][0] = 1292ns;
slave_timing[1][5].t_rxd2[1][2] = 2016ns;
slave_timing[1][5].t_rxd2[2][1] = 1688ns;

slave_timing[1][6].info_corner          = 0;
slave_timing[1][6].info_temp__j__       = 25;
slave_timing[1][6].info_i__quite_rec__  = 0.006000000;
slave_timing[1][6].info_dtr__ib__       = 1;
slave_timing[1][6].info_i__offset_rec__ = -0.001000000;
slave_timing[1][6].info_i__max_slave__  = 0.027000000;
slave_timing[1][6].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][6].info_r__dsi_bus__    = 5.000;

slave_timing[1][6].t_rxd1[0][1] = 1879ns;
slave_timing[1][6].t_rxd1[1][0] = 1682ns;
slave_timing[1][6].t_rxd1[0][2] = 1375ns;
slave_timing[1][6].t_rxd1[2][0] = 2049ns;
slave_timing[1][6].t_rxd2[0][2] = 2012ns;
slave_timing[1][6].t_rxd2[2][0] = 1413ns;
slave_timing[1][6].t_rxd2[1][2] = 1634ns;
slave_timing[1][6].t_rxd2[2][1] = 1954ns;

slave_timing[1][7].info_corner          = 0;
slave_timing[1][7].info_temp__j__       = 25;
slave_timing[1][7].info_i__quite_rec__  = 0.006000000;
slave_timing[1][7].info_dtr__ib__       = 1;
slave_timing[1][7].info_i__offset_rec__ = 0.001000000;
slave_timing[1][7].info_i__max_slave__  = 0.027000000;
slave_timing[1][7].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][7].info_r__dsi_bus__    = 5.000;

slave_timing[1][7].t_rxd1[0][1] = 1678ns;
slave_timing[1][7].t_rxd1[1][0] = 1882ns;
slave_timing[1][7].t_rxd1[0][2] = 1265ns;
slave_timing[1][7].t_rxd1[2][0] = 2205ns;
slave_timing[1][7].t_rxd2[0][2] = 1879ns;
slave_timing[1][7].t_rxd2[2][0] = 1508ns;
slave_timing[1][7].t_rxd2[1][2] = 1446ns;
slave_timing[1][7].t_rxd2[2][1] = 2250ns;

slave_timing[1][8].info_corner          = 0;
slave_timing[1][8].info_temp__j__       = 25;
slave_timing[1][8].info_i__quite_rec__  = 0.006000000;
slave_timing[1][8].info_dtr__ib__       = -1;
slave_timing[1][8].info_i__offset_rec__ = -0.001000000;
slave_timing[1][8].info_i__max_slave__  = 0.021000000;
slave_timing[1][8].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][8].info_r__dsi_bus__    = 5.000;

slave_timing[1][8].t_rxd1[0][1] = 2431ns;
slave_timing[1][8].t_rxd1[1][0] = 1751ns;
slave_timing[1][8].t_rxd1[0][2] = 1679ns;
slave_timing[1][8].t_rxd1[2][0] = 2205ns;
slave_timing[1][8].t_rxd2[0][2] = 2755ns;
slave_timing[1][8].t_rxd2[2][0] = 1388ns;
slave_timing[1][8].t_rxd2[1][2] = 2455ns;
slave_timing[1][8].t_rxd2[2][1] = 1755ns;

slave_timing[1][9].info_corner          = 0;
slave_timing[1][9].info_temp__j__       = 25;
slave_timing[1][9].info_i__quite_rec__  = 0.006000000;
slave_timing[1][9].info_dtr__ib__       = -1;
slave_timing[1][9].info_i__offset_rec__ = 0.001000000;
slave_timing[1][9].info_i__max_slave__  = 0.021000000;
slave_timing[1][9].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][9].info_r__dsi_bus__    = 5.000;

slave_timing[1][9].t_rxd1[0][1] = 2039ns;
slave_timing[1][9].t_rxd1[1][0] = 2049ns;
slave_timing[1][9].t_rxd1[0][2] = 1532ns;
slave_timing[1][9].t_rxd1[2][0] = 2429ns;
slave_timing[1][9].t_rxd2[0][2] = 2421ns;
slave_timing[1][9].t_rxd2[2][0] = 1548ns;
slave_timing[1][9].t_rxd2[1][2] = 2057ns;
slave_timing[1][9].t_rxd2[2][1] = 2055ns;

slave_timing[1][10].info_corner          = 0;
slave_timing[1][10].info_temp__j__       = 25;
slave_timing[1][10].info_i__quite_rec__  = 0.006000000;
slave_timing[1][10].info_dtr__ib__       = -1;
slave_timing[1][10].info_i__offset_rec__ = -0.001000000;
slave_timing[1][10].info_i__max_slave__  = 0.027000000;
slave_timing[1][10].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][10].info_r__dsi_bus__    = 5.000;

slave_timing[1][10].t_rxd1[0][1] = 2053ns;
slave_timing[1][10].t_rxd1[1][0] = 1933ns;
slave_timing[1][10].t_rxd1[0][2] = 1535ns;
slave_timing[1][10].t_rxd1[2][0] = 2333ns;
slave_timing[1][10].t_rxd2[0][2] = 2174ns;
slave_timing[1][10].t_rxd2[2][0] = 1661ns;
slave_timing[1][10].t_rxd2[1][2] = 1712ns;
slave_timing[1][10].t_rxd2[2][1] = 2361ns;

slave_timing[1][11].info_corner          = 0;
slave_timing[1][11].info_temp__j__       = 25;
slave_timing[1][11].info_i__quite_rec__  = 0.006000000;
slave_timing[1][11].info_dtr__ib__       = -1;
slave_timing[1][11].info_i__offset_rec__ = 0.001000000;
slave_timing[1][11].info_i__max_slave__  = 0.027000000;
slave_timing[1][11].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][11].info_r__dsi_bus__    = 5.000;

slave_timing[1][11].t_rxd1[0][1] = 1813ns;
slave_timing[1][11].t_rxd1[1][0] = 2192ns;
slave_timing[1][11].t_rxd1[0][2] = 1410ns;
slave_timing[1][11].t_rxd1[2][0] = 2543ns;
slave_timing[1][11].t_rxd2[0][2] = 2037ns;
slave_timing[1][11].t_rxd2[2][0] = 1773ns;
slave_timing[1][11].t_rxd2[1][2] = 1479ns;
slave_timing[1][11].t_rxd2[2][1] = 2962ns;

slave_timing[1][12].info_corner          = 0;
slave_timing[1][12].info_temp__j__       = 25;
slave_timing[1][12].info_i__quite_rec__  = 0.006000000;
slave_timing[1][12].info_dtr__ib__       = 1;
slave_timing[1][12].info_i__offset_rec__ = -0.001000000;
slave_timing[1][12].info_i__max_slave__  = 0.021000000;
slave_timing[1][12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][12].info_r__dsi_bus__    = 5.000;

slave_timing[1][12].t_rxd1[0][1] = 2564ns;
slave_timing[1][12].t_rxd1[1][0] = 1706ns;
slave_timing[1][12].t_rxd1[0][2] = 1714ns;
slave_timing[1][12].t_rxd1[2][0] = 2177ns;
slave_timing[1][12].t_rxd2[0][2] = 3143ns;
slave_timing[1][12].t_rxd2[2][0] = 1297ns;
slave_timing[1][12].t_rxd2[1][2] = 2878ns;
slave_timing[1][12].t_rxd2[2][1] = 1614ns;

slave_timing[1][13].info_corner          = 0;
slave_timing[1][13].info_temp__j__       = 25;
slave_timing[1][13].info_i__quite_rec__  = 0.006000000;
slave_timing[1][13].info_dtr__ib__       = 1;
slave_timing[1][13].info_i__offset_rec__ = 0.001000000;
slave_timing[1][13].info_i__max_slave__  = 0.021000000;
slave_timing[1][13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][13].info_r__dsi_bus__    = 5.000;

slave_timing[1][13].t_rxd1[0][1] = 2118ns;
slave_timing[1][13].t_rxd1[1][0] = 2004ns;
slave_timing[1][13].t_rxd1[0][2] = 1566ns;
slave_timing[1][13].t_rxd1[2][0] = 2390ns;
slave_timing[1][13].t_rxd2[0][2] = 2590ns;
slave_timing[1][13].t_rxd2[2][0] = 1470ns;
slave_timing[1][13].t_rxd2[1][2] = 2265ns;
slave_timing[1][13].t_rxd2[2][1] = 1905ns;

slave_timing[1][14].info_corner          = 0;
slave_timing[1][14].info_temp__j__       = 25;
slave_timing[1][14].info_i__quite_rec__  = 0.006000000;
slave_timing[1][14].info_dtr__ib__       = 1;
slave_timing[1][14].info_i__offset_rec__ = -0.001000000;
slave_timing[1][14].info_i__max_slave__  = 0.027000000;
slave_timing[1][14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][14].info_r__dsi_bus__    = 5.000;

slave_timing[1][14].t_rxd1[0][1] = 2116ns;
slave_timing[1][14].t_rxd1[1][0] = 1900ns;
slave_timing[1][14].t_rxd1[0][2] = 1562ns;
slave_timing[1][14].t_rxd1[2][0] = 2307ns;
slave_timing[1][14].t_rxd2[0][2] = 2261ns;
slave_timing[1][14].t_rxd2[2][0] = 1604ns;
slave_timing[1][14].t_rxd2[1][2] = 1845ns;
slave_timing[1][14].t_rxd2[2][1] = 2198ns;

slave_timing[1][15].info_corner          = 0;
slave_timing[1][15].info_temp__j__       = 25;
slave_timing[1][15].info_i__quite_rec__  = 0.006000000;
slave_timing[1][15].info_dtr__ib__       = 1;
slave_timing[1][15].info_i__offset_rec__ = 0.001000000;
slave_timing[1][15].info_i__max_slave__  = 0.027000000;
slave_timing[1][15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][15].info_r__dsi_bus__    = 5.000;

slave_timing[1][15].t_rxd1[0][1] = 1890ns;
slave_timing[1][15].t_rxd1[1][0] = 2121ns;
slave_timing[1][15].t_rxd1[0][2] = 1440ns;
slave_timing[1][15].t_rxd1[2][0] = 2483ns;
slave_timing[1][15].t_rxd2[0][2] = 2114ns;
slave_timing[1][15].t_rxd2[2][0] = 1706ns;
slave_timing[1][15].t_rxd2[1][2] = 1636ns;
slave_timing[1][15].t_rxd2[2][1] = 2535ns;

slave_timing[1][16].info_corner          = 0;
slave_timing[1][16].info_temp__j__       = 25;
slave_timing[1][16].info_i__quite_rec__  = 0.003000000;
slave_timing[1][16].info_dtr__ib__       = -1;
slave_timing[1][16].info_i__offset_rec__ = -0.001000000;
slave_timing[1][16].info_i__max_slave__  = 0.021000000;
slave_timing[1][16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][16].info_r__dsi_bus__    = 5.000;

slave_timing[1][16].t_rxd1[0][1] = 2146ns;
slave_timing[1][16].t_rxd1[1][0] = 1558ns;
slave_timing[1][16].t_rxd1[0][2] = 1478ns;
slave_timing[1][16].t_rxd1[2][0] = 1966ns;
slave_timing[1][16].t_rxd2[0][2] = 2433ns;
slave_timing[1][16].t_rxd2[2][0] = 1221ns;
slave_timing[1][16].t_rxd2[1][2] = 2170ns;
slave_timing[1][16].t_rxd2[2][1] = 1561ns;

slave_timing[1][17].info_corner          = 0;
slave_timing[1][17].info_temp__j__       = 25;
slave_timing[1][17].info_i__quite_rec__  = 0.003000000;
slave_timing[1][17].info_dtr__ib__       = -1;
slave_timing[1][17].info_i__offset_rec__ = 0.001000000;
slave_timing[1][17].info_i__max_slave__  = 0.021000000;
slave_timing[1][17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][17].info_r__dsi_bus__    = 5.000;

slave_timing[1][17].t_rxd1[0][1] = 1799ns;
slave_timing[1][17].t_rxd1[1][0] = 1833ns;
slave_timing[1][17].t_rxd1[0][2] = 1343ns;
slave_timing[1][17].t_rxd1[2][0] = 2163ns;
slave_timing[1][17].t_rxd2[0][2] = 2143ns;
slave_timing[1][17].t_rxd2[2][0] = 1367ns;
slave_timing[1][17].t_rxd2[1][2] = 1813ns;
slave_timing[1][17].t_rxd2[2][1] = 1839ns;

slave_timing[1][18].info_corner          = 0;
slave_timing[1][18].info_temp__j__       = 25;
slave_timing[1][18].info_i__quite_rec__  = 0.003000000;
slave_timing[1][18].info_dtr__ib__       = -1;
slave_timing[1][18].info_i__offset_rec__ = -0.001000000;
slave_timing[1][18].info_i__max_slave__  = 0.027000000;
slave_timing[1][18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][18].info_r__dsi_bus__    = 5.000;

slave_timing[1][18].t_rxd1[0][1] = 1816ns;
slave_timing[1][18].t_rxd1[1][0] = 1720ns;
slave_timing[1][18].t_rxd1[0][2] = 1357ns;
slave_timing[1][18].t_rxd1[2][0] = 2063ns;
slave_timing[1][18].t_rxd2[0][2] = 1938ns;
slave_timing[1][18].t_rxd2[2][0] = 1461ns;
slave_timing[1][18].t_rxd2[1][2] = 1504ns;
slave_timing[1][18].t_rxd2[2][1] = 2107ns;

slave_timing[1][19].info_corner          = 0;
slave_timing[1][19].info_temp__j__       = 25;
slave_timing[1][19].info_i__quite_rec__  = 0.003000000;
slave_timing[1][19].info_dtr__ib__       = -1;
slave_timing[1][19].info_i__offset_rec__ = 0.001000000;
slave_timing[1][19].info_i__max_slave__  = 0.027000000;
slave_timing[1][19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][19].info_r__dsi_bus__    = 5.000;

slave_timing[1][19].t_rxd1[0][1] = 1598ns;
slave_timing[1][19].t_rxd1[1][0] = 1955ns;
slave_timing[1][19].t_rxd1[0][2] = 1233ns;
slave_timing[1][19].t_rxd1[2][0] = 2263ns;
slave_timing[1][19].t_rxd2[0][2] = 1804ns;
slave_timing[1][19].t_rxd2[2][0] = 1574ns;
slave_timing[1][19].t_rxd2[1][2] = 1292ns;
slave_timing[1][19].t_rxd2[2][1] = 2666ns;

slave_timing[1][20].info_corner          = 0;
slave_timing[1][20].info_temp__j__       = 25;
slave_timing[1][20].info_i__quite_rec__  = 0.003000000;
slave_timing[1][20].info_dtr__ib__       = 1;
slave_timing[1][20].info_i__offset_rec__ = -0.001000000;
slave_timing[1][20].info_i__max_slave__  = 0.021000000;
slave_timing[1][20].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][20].info_r__dsi_bus__    = 5.000;

slave_timing[1][20].t_rxd1[0][1] = 2262ns;
slave_timing[1][20].t_rxd1[1][0] = 1519ns;
slave_timing[1][20].t_rxd1[0][2] = 1509ns;
slave_timing[1][20].t_rxd1[2][0] = 1941ns;
slave_timing[1][20].t_rxd2[0][2] = 2763ns;
slave_timing[1][20].t_rxd2[2][0] = 1140ns;
slave_timing[1][20].t_rxd2[1][2] = 2529ns;
slave_timing[1][20].t_rxd2[2][1] = 1432ns;

slave_timing[1][21].info_corner          = 0;
slave_timing[1][21].info_temp__j__       = 25;
slave_timing[1][21].info_i__quite_rec__  = 0.003000000;
slave_timing[1][21].info_dtr__ib__       = 1;
slave_timing[1][21].info_i__offset_rec__ = 0.001000000;
slave_timing[1][21].info_i__max_slave__  = 0.021000000;
slave_timing[1][21].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][21].info_r__dsi_bus__    = 5.000;

slave_timing[1][21].t_rxd1[0][1] = 1871ns;
slave_timing[1][21].t_rxd1[1][0] = 1791ns;
slave_timing[1][21].t_rxd1[0][2] = 1373ns;
slave_timing[1][21].t_rxd1[2][0] = 2130ns;
slave_timing[1][21].t_rxd2[0][2] = 2290ns;
slave_timing[1][21].t_rxd2[2][0] = 1297ns;
slave_timing[1][21].t_rxd2[1][2] = 2002ns;
slave_timing[1][21].t_rxd2[2][1] = 1698ns;

slave_timing[1][22].info_corner          = 0;
slave_timing[1][22].info_temp__j__       = 25;
slave_timing[1][22].info_i__quite_rec__  = 0.003000000;
slave_timing[1][22].info_dtr__ib__       = 1;
slave_timing[1][22].info_i__offset_rec__ = -0.001000000;
slave_timing[1][22].info_i__max_slave__  = 0.027000000;
slave_timing[1][22].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][22].info_r__dsi_bus__    = 5.000;

slave_timing[1][22].t_rxd1[0][1] = 1873ns;
slave_timing[1][22].t_rxd1[1][0] = 1687ns;
slave_timing[1][22].t_rxd1[0][2] = 1373ns;
slave_timing[1][22].t_rxd1[2][0] = 2053ns;
slave_timing[1][22].t_rxd2[0][2] = 2006ns;
slave_timing[1][22].t_rxd2[2][0] = 1417ns;
slave_timing[1][22].t_rxd2[1][2] = 1622ns;
slave_timing[1][22].t_rxd2[2][1] = 1964ns;

slave_timing[1][23].info_corner          = 0;
slave_timing[1][23].info_temp__j__       = 25;
slave_timing[1][23].info_i__quite_rec__  = 0.003000000;
slave_timing[1][23].info_dtr__ib__       = 1;
slave_timing[1][23].info_i__offset_rec__ = 0.001000000;
slave_timing[1][23].info_i__max_slave__  = 0.027000000;
slave_timing[1][23].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][23].info_r__dsi_bus__    = 5.000;

slave_timing[1][23].t_rxd1[0][1] = 1670ns;
slave_timing[1][23].t_rxd1[1][0] = 1892ns;
slave_timing[1][23].t_rxd1[0][2] = 1274ns;
slave_timing[1][23].t_rxd1[2][0] = 2208ns;
slave_timing[1][23].t_rxd2[0][2] = 1884ns;
slave_timing[1][23].t_rxd2[2][0] = 1512ns;
slave_timing[1][23].t_rxd2[1][2] = 1439ns;
slave_timing[1][23].t_rxd2[2][1] = 2264ns;

slave_timing[1][24].info_corner          = 0;
slave_timing[1][24].info_temp__j__       = 25;
slave_timing[1][24].info_i__quite_rec__  = 0.003000000;
slave_timing[1][24].info_dtr__ib__       = -1;
slave_timing[1][24].info_i__offset_rec__ = -0.001000000;
slave_timing[1][24].info_i__max_slave__  = 0.021000000;
slave_timing[1][24].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][24].info_r__dsi_bus__    = 5.000;

slave_timing[1][24].t_rxd1[0][1] = 2409ns;
slave_timing[1][24].t_rxd1[1][0] = 1761ns;
slave_timing[1][24].t_rxd1[0][2] = 1674ns;
slave_timing[1][24].t_rxd1[2][0] = 2210ns;
slave_timing[1][24].t_rxd2[0][2] = 2735ns;
slave_timing[1][24].t_rxd2[2][0] = 1394ns;
slave_timing[1][24].t_rxd2[1][2] = 2433ns;
slave_timing[1][24].t_rxd2[2][1] = 1767ns;

slave_timing[1][25].info_corner          = 0;
slave_timing[1][25].info_temp__j__       = 25;
slave_timing[1][25].info_i__quite_rec__  = 0.003000000;
slave_timing[1][25].info_dtr__ib__       = -1;
slave_timing[1][25].info_i__offset_rec__ = 0.001000000;
slave_timing[1][25].info_i__max_slave__  = 0.021000000;
slave_timing[1][25].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][25].info_r__dsi_bus__    = 5.000;

slave_timing[1][25].t_rxd1[0][1] = 2024ns;
slave_timing[1][25].t_rxd1[1][0] = 2060ns;
slave_timing[1][25].t_rxd1[0][2] = 1525ns;
slave_timing[1][25].t_rxd1[2][0] = 2435ns;
slave_timing[1][25].t_rxd2[0][2] = 2408ns;
slave_timing[1][25].t_rxd2[2][0] = 1552ns;
slave_timing[1][25].t_rxd2[1][2] = 2039ns;
slave_timing[1][25].t_rxd2[2][1] = 2068ns;

slave_timing[1][26].info_corner          = 0;
slave_timing[1][26].info_temp__j__       = 25;
slave_timing[1][26].info_i__quite_rec__  = 0.003000000;
slave_timing[1][26].info_dtr__ib__       = -1;
slave_timing[1][26].info_i__offset_rec__ = -0.001000000;
slave_timing[1][26].info_i__max_slave__  = 0.027000000;
slave_timing[1][26].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][26].info_r__dsi_bus__    = 5.000;

slave_timing[1][26].t_rxd1[0][1] = 2042ns;
slave_timing[1][26].t_rxd1[1][0] = 1941ns;
slave_timing[1][26].t_rxd1[0][2] = 1532ns;
slave_timing[1][26].t_rxd1[2][0] = 2338ns;
slave_timing[1][26].t_rxd2[0][2] = 2167ns;
slave_timing[1][26].t_rxd2[2][0] = 1665ns;
slave_timing[1][26].t_rxd2[1][2] = 1702ns;
slave_timing[1][26].t_rxd2[2][1] = 2372ns;

slave_timing[1][27].info_corner          = 0;
slave_timing[1][27].info_temp__j__       = 25;
slave_timing[1][27].info_i__quite_rec__  = 0.003000000;
slave_timing[1][27].info_dtr__ib__       = -1;
slave_timing[1][27].info_i__offset_rec__ = 0.001000000;
slave_timing[1][27].info_i__max_slave__  = 0.027000000;
slave_timing[1][27].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][27].info_r__dsi_bus__    = 5.000;

slave_timing[1][27].t_rxd1[0][1] = 1802ns;
slave_timing[1][27].t_rxd1[1][0] = 2201ns;
slave_timing[1][27].t_rxd1[0][2] = 1408ns;
slave_timing[1][27].t_rxd1[2][0] = 2550ns;
slave_timing[1][27].t_rxd2[0][2] = 2032ns;
slave_timing[1][27].t_rxd2[2][0] = 1779ns;
slave_timing[1][27].t_rxd2[1][2] = 1469ns;
slave_timing[1][27].t_rxd2[2][1] = 3004ns;

slave_timing[1][28].info_corner          = 0;
slave_timing[1][28].info_temp__j__       = 25;
slave_timing[1][28].info_i__quite_rec__  = 0.003000000;
slave_timing[1][28].info_dtr__ib__       = 1;
slave_timing[1][28].info_i__offset_rec__ = -0.001000000;
slave_timing[1][28].info_i__max_slave__  = 0.021000000;
slave_timing[1][28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][28].info_r__dsi_bus__    = 5.000;

slave_timing[1][28].t_rxd1[0][1] = 2537ns;
slave_timing[1][28].t_rxd1[1][0] = 1717ns;
slave_timing[1][28].t_rxd1[0][2] = 1709ns;
slave_timing[1][28].t_rxd1[2][0] = 2182ns;
slave_timing[1][28].t_rxd2[0][2] = 3106ns;
slave_timing[1][28].t_rxd2[2][0] = 1303ns;
slave_timing[1][28].t_rxd2[1][2] = 2836ns;
slave_timing[1][28].t_rxd2[2][1] = 1624ns;

slave_timing[1][29].info_corner          = 0;
slave_timing[1][29].info_temp__j__       = 25;
slave_timing[1][29].info_i__quite_rec__  = 0.003000000;
slave_timing[1][29].info_dtr__ib__       = 1;
slave_timing[1][29].info_i__offset_rec__ = 0.001000000;
slave_timing[1][29].info_i__max_slave__  = 0.021000000;
slave_timing[1][29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][29].info_r__dsi_bus__    = 5.000;

slave_timing[1][29].t_rxd1[0][1] = 2103ns;
slave_timing[1][29].t_rxd1[1][0] = 2014ns;
slave_timing[1][29].t_rxd1[0][2] = 1561ns;
slave_timing[1][29].t_rxd1[2][0] = 2397ns;
slave_timing[1][29].t_rxd2[0][2] = 2576ns;
slave_timing[1][29].t_rxd2[2][0] = 1477ns;
slave_timing[1][29].t_rxd2[1][2] = 2250ns;
slave_timing[1][29].t_rxd2[2][1] = 1915ns;

slave_timing[1][30].info_corner          = 0;
slave_timing[1][30].info_temp__j__       = 25;
slave_timing[1][30].info_i__quite_rec__  = 0.003000000;
slave_timing[1][30].info_dtr__ib__       = 1;
slave_timing[1][30].info_i__offset_rec__ = -0.001000000;
slave_timing[1][30].info_i__max_slave__  = 0.027000000;
slave_timing[1][30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][30].info_r__dsi_bus__    = 5.000;

slave_timing[1][30].t_rxd1[0][1] = 2103ns;
slave_timing[1][30].t_rxd1[1][0] = 1903ns;
slave_timing[1][30].t_rxd1[0][2] = 1559ns;
slave_timing[1][30].t_rxd1[2][0] = 2310ns;
slave_timing[1][30].t_rxd2[0][2] = 2254ns;
slave_timing[1][30].t_rxd2[2][0] = 1609ns;
slave_timing[1][30].t_rxd2[1][2] = 1835ns;
slave_timing[1][30].t_rxd2[2][1] = 2207ns;

slave_timing[1][31].info_corner          = 0;
slave_timing[1][31].info_temp__j__       = 25;
slave_timing[1][31].info_i__quite_rec__  = 0.003000000;
slave_timing[1][31].info_dtr__ib__       = 1;
slave_timing[1][31].info_i__offset_rec__ = 0.001000000;
slave_timing[1][31].info_i__max_slave__  = 0.027000000;
slave_timing[1][31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][31].info_r__dsi_bus__    = 5.000;

slave_timing[1][31].t_rxd1[0][1] = 1881ns;
slave_timing[1][31].t_rxd1[1][0] = 2128ns;
slave_timing[1][31].t_rxd1[0][2] = 1450ns;
slave_timing[1][31].t_rxd1[2][0] = 2488ns;
slave_timing[1][31].t_rxd2[0][2] = 2121ns;
slave_timing[1][31].t_rxd2[2][0] = 1710ns;
slave_timing[1][31].t_rxd2[1][2] = 1631ns;
slave_timing[1][31].t_rxd2[2][1] = 2548ns;

slave_timing[1][32].info_corner          = 0;
slave_timing[1][32].info_temp__j__       = 25;
slave_timing[1][32].info_i__quite_rec__  = 0.000000000;
slave_timing[1][32].info_dtr__ib__       = -1;
slave_timing[1][32].info_i__offset_rec__ = -0.001000000;
slave_timing[1][32].info_i__max_slave__  = 0.021000000;
slave_timing[1][32].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][32].info_r__dsi_bus__    = 5.000;

slave_timing[1][32].t_rxd1[0][1] = 2171ns;
slave_timing[1][32].t_rxd1[1][0] = 1549ns;
slave_timing[1][32].t_rxd1[0][2] = 1483ns;
slave_timing[1][32].t_rxd1[2][0] = 1961ns;
slave_timing[1][32].t_rxd2[0][2] = 2453ns;
slave_timing[1][32].t_rxd2[2][0] = 1215ns;
slave_timing[1][32].t_rxd2[1][2] = 2193ns;
slave_timing[1][32].t_rxd2[2][1] = 1553ns;

slave_timing[1][33].info_corner          = 0;
slave_timing[1][33].info_temp__j__       = 25;
slave_timing[1][33].info_i__quite_rec__  = 0.000000000;
slave_timing[1][33].info_dtr__ib__       = -1;
slave_timing[1][33].info_i__offset_rec__ = 0.001000000;
slave_timing[1][33].info_i__max_slave__  = 0.021000000;
slave_timing[1][33].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][33].info_r__dsi_bus__    = 5.000;

slave_timing[1][33].t_rxd1[0][1] = 1816ns;
slave_timing[1][33].t_rxd1[1][0] = 1823ns;
slave_timing[1][33].t_rxd1[0][2] = 1348ns;
slave_timing[1][33].t_rxd1[2][0] = 2155ns;
slave_timing[1][33].t_rxd2[0][2] = 2156ns;
slave_timing[1][33].t_rxd2[2][0] = 1360ns;
slave_timing[1][33].t_rxd2[1][2] = 1829ns;
slave_timing[1][33].t_rxd2[2][1] = 1827ns;

slave_timing[1][34].info_corner          = 0;
slave_timing[1][34].info_temp__j__       = 25;
slave_timing[1][34].info_i__quite_rec__  = 0.000000000;
slave_timing[1][34].info_dtr__ib__       = -1;
slave_timing[1][34].info_i__offset_rec__ = -0.001000000;
slave_timing[1][34].info_i__max_slave__  = 0.027000000;
slave_timing[1][34].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][34].info_r__dsi_bus__    = 5.000;

slave_timing[1][34].t_rxd1[0][1] = 1826ns;
slave_timing[1][34].t_rxd1[1][0] = 1713ns;
slave_timing[1][34].t_rxd1[0][2] = 1362ns;
slave_timing[1][34].t_rxd1[2][0] = 2057ns;
slave_timing[1][34].t_rxd2[0][2] = 1946ns;
slave_timing[1][34].t_rxd2[2][0] = 1454ns;
slave_timing[1][34].t_rxd2[1][2] = 1514ns;
slave_timing[1][34].t_rxd2[2][1] = 2094ns;

slave_timing[1][35].info_corner          = 0;
slave_timing[1][35].info_temp__j__       = 25;
slave_timing[1][35].info_i__quite_rec__  = 0.000000000;
slave_timing[1][35].info_dtr__ib__       = -1;
slave_timing[1][35].info_i__offset_rec__ = 0.001000000;
slave_timing[1][35].info_i__max_slave__  = 0.027000000;
slave_timing[1][35].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][35].info_r__dsi_bus__    = 5.000;

slave_timing[1][35].t_rxd1[0][1] = 1607ns;
slave_timing[1][35].t_rxd1[1][0] = 1947ns;
slave_timing[1][35].t_rxd1[0][2] = 1236ns;
slave_timing[1][35].t_rxd1[2][0] = 2255ns;
slave_timing[1][35].t_rxd2[0][2] = 1811ns;
slave_timing[1][35].t_rxd2[2][0] = 1569ns;
slave_timing[1][35].t_rxd2[1][2] = 1302ns;
slave_timing[1][35].t_rxd2[2][1] = 2621ns;

slave_timing[1][36].info_corner          = 0;
slave_timing[1][36].info_temp__j__       = 25;
slave_timing[1][36].info_i__quite_rec__  = 0.000000000;
slave_timing[1][36].info_dtr__ib__       = 1;
slave_timing[1][36].info_i__offset_rec__ = -0.001000000;
slave_timing[1][36].info_i__max_slave__  = 0.021000000;
slave_timing[1][36].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][36].info_r__dsi_bus__    = 5.000;

slave_timing[1][36].t_rxd1[0][1] = 2357ns;
slave_timing[1][36].t_rxd1[1][0] = 1475ns;
slave_timing[1][36].t_rxd1[0][2] = 1531ns;
slave_timing[1][36].t_rxd1[2][0] = 1917ns;
slave_timing[1][36].t_rxd2[0][2] = 2936ns;
slave_timing[1][36].t_rxd2[2][0] = 1111ns;
slave_timing[1][36].t_rxd2[1][2] = 2706ns;
slave_timing[1][36].t_rxd2[2][1] = 1388ns;

slave_timing[1][37].info_corner          = 0;
slave_timing[1][37].info_temp__j__       = 25;
slave_timing[1][37].info_i__quite_rec__  = 0.000000000;
slave_timing[1][37].info_dtr__ib__       = 1;
slave_timing[1][37].info_i__offset_rec__ = 0.001000000;
slave_timing[1][37].info_i__max_slave__  = 0.021000000;
slave_timing[1][37].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][37].info_r__dsi_bus__    = 5.000;

slave_timing[1][37].t_rxd1[0][1] = 1924ns;
slave_timing[1][37].t_rxd1[1][0] = 1746ns;
slave_timing[1][37].t_rxd1[0][2] = 1395ns;
slave_timing[1][37].t_rxd1[2][0] = 2097ns;
slave_timing[1][37].t_rxd2[0][2] = 2341ns;
slave_timing[1][37].t_rxd2[2][0] = 1275ns;
slave_timing[1][37].t_rxd2[1][2] = 2061ns;
slave_timing[1][37].t_rxd2[2][1] = 1657ns;

slave_timing[1][38].info_corner          = 0;
slave_timing[1][38].info_temp__j__       = 25;
slave_timing[1][38].info_i__quite_rec__  = 0.000000000;
slave_timing[1][38].info_dtr__ib__       = 1;
slave_timing[1][38].info_i__offset_rec__ = -0.001000000;
slave_timing[1][38].info_i__max_slave__  = 0.027000000;
slave_timing[1][38].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][38].info_r__dsi_bus__    = 5.000;

slave_timing[1][38].t_rxd1[0][1] = 1887ns;
slave_timing[1][38].t_rxd1[1][0] = 1677ns;
slave_timing[1][38].t_rxd1[0][2] = 1378ns;
slave_timing[1][38].t_rxd1[2][0] = 2046ns;
slave_timing[1][38].t_rxd2[0][2] = 2015ns;
slave_timing[1][38].t_rxd2[2][0] = 1410ns;
slave_timing[1][38].t_rxd2[1][2] = 1638ns;
slave_timing[1][38].t_rxd2[2][1] = 1947ns;

slave_timing[1][39].info_corner          = 0;
slave_timing[1][39].info_temp__j__       = 25;
slave_timing[1][39].info_i__quite_rec__  = 0.000000000;
slave_timing[1][39].info_dtr__ib__       = 1;
slave_timing[1][39].info_i__offset_rec__ = 0.001000000;
slave_timing[1][39].info_i__max_slave__  = 0.027000000;
slave_timing[1][39].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][39].info_r__dsi_bus__    = 5.000;

slave_timing[1][39].t_rxd1[0][1] = 1659ns;
slave_timing[1][39].t_rxd1[1][0] = 1904ns;
slave_timing[1][39].t_rxd1[0][2] = 1267ns;
slave_timing[1][39].t_rxd1[2][0] = 2220ns;
slave_timing[1][39].t_rxd2[0][2] = 1882ns;
slave_timing[1][39].t_rxd2[2][0] = 1515ns;
slave_timing[1][39].t_rxd2[1][2] = 1431ns;
slave_timing[1][39].t_rxd2[2][1] = 2277ns;

slave_timing[1][40].info_corner          = 0;
slave_timing[1][40].info_temp__j__       = 25;
slave_timing[1][40].info_i__quite_rec__  = 0.000000000;
slave_timing[1][40].info_dtr__ib__       = -1;
slave_timing[1][40].info_i__offset_rec__ = -0.001000000;
slave_timing[1][40].info_i__max_slave__  = 0.021000000;
slave_timing[1][40].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][40].info_r__dsi_bus__    = 5.000;

slave_timing[1][40].t_rxd1[0][1] = 2487ns;
slave_timing[1][40].t_rxd1[1][0] = 1723ns;
slave_timing[1][40].t_rxd1[0][2] = 1695ns;
slave_timing[1][40].t_rxd1[2][0] = 2186ns;
slave_timing[1][40].t_rxd2[0][2] = 2806ns;
slave_timing[1][40].t_rxd2[2][0] = 1370ns;
slave_timing[1][40].t_rxd2[1][2] = 2514ns;
slave_timing[1][40].t_rxd2[2][1] = 1726ns;

slave_timing[1][41].info_corner          = 0;
slave_timing[1][41].info_temp__j__       = 25;
slave_timing[1][41].info_i__quite_rec__  = 0.000000000;
slave_timing[1][41].info_dtr__ib__       = -1;
slave_timing[1][41].info_i__offset_rec__ = 0.001000000;
slave_timing[1][41].info_i__max_slave__  = 0.021000000;
slave_timing[1][41].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][41].info_r__dsi_bus__    = 5.000;

slave_timing[1][41].t_rxd1[0][1] = 2073ns;
slave_timing[1][41].t_rxd1[1][0] = 2019ns;
slave_timing[1][41].t_rxd1[0][2] = 1547ns;
slave_timing[1][41].t_rxd1[2][0] = 2400ns;
slave_timing[1][41].t_rxd2[0][2] = 2447ns;
slave_timing[1][41].t_rxd2[2][0] = 1531ns;
slave_timing[1][41].t_rxd2[1][2] = 2091ns;
slave_timing[1][41].t_rxd2[2][1] = 2024ns;

slave_timing[1][42].info_corner          = 0;
slave_timing[1][42].info_temp__j__       = 25;
slave_timing[1][42].info_i__quite_rec__  = 0.000000000;
slave_timing[1][42].info_dtr__ib__       = -1;
slave_timing[1][42].info_i__offset_rec__ = -0.001000000;
slave_timing[1][42].info_i__max_slave__  = 0.027000000;
slave_timing[1][42].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][42].info_r__dsi_bus__    = 5.000;

slave_timing[1][42].t_rxd1[0][1] = 2080ns;
slave_timing[1][42].t_rxd1[1][0] = 1908ns;
slave_timing[1][42].t_rxd1[0][2] = 1548ns;
slave_timing[1][42].t_rxd1[2][0] = 2315ns;
slave_timing[1][42].t_rxd2[0][2] = 2190ns;
slave_timing[1][42].t_rxd2[2][0] = 1651ns;
slave_timing[1][42].t_rxd2[1][2] = 1736ns;
slave_timing[1][42].t_rxd2[2][1] = 2322ns;

slave_timing[1][43].info_corner          = 0;
slave_timing[1][43].info_temp__j__       = 25;
slave_timing[1][43].info_i__quite_rec__  = 0.000000000;
slave_timing[1][43].info_dtr__ib__       = -1;
slave_timing[1][43].info_i__offset_rec__ = 0.001000000;
slave_timing[1][43].info_i__max_slave__  = 0.027000000;
slave_timing[1][43].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][43].info_r__dsi_bus__    = 5.000;

slave_timing[1][43].t_rxd1[0][1] = 1838ns;
slave_timing[1][43].t_rxd1[1][0] = 2161ns;
slave_timing[1][43].t_rxd1[0][2] = 1426ns;
slave_timing[1][43].t_rxd1[2][0] = 2517ns;
slave_timing[1][43].t_rxd2[0][2] = 2052ns;
slave_timing[1][43].t_rxd2[2][0] = 1763ns;
slave_timing[1][43].t_rxd2[1][2] = 1506ns;
slave_timing[1][43].t_rxd2[2][1] = 2853ns;

slave_timing[1][44].info_corner          = 0;
slave_timing[1][44].info_temp__j__       = 25;
slave_timing[1][44].info_i__quite_rec__  = 0.000000000;
slave_timing[1][44].info_dtr__ib__       = 1;
slave_timing[1][44].info_i__offset_rec__ = -0.001000000;
slave_timing[1][44].info_i__max_slave__  = 0.021000000;
slave_timing[1][44].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][44].info_r__dsi_bus__    = 5.000;

slave_timing[1][44].t_rxd1[0][1] = 2576ns;
slave_timing[1][44].t_rxd1[1][0] = 1703ns;
slave_timing[1][44].t_rxd1[0][2] = 1733ns;
slave_timing[1][44].t_rxd1[2][0] = 2154ns;
slave_timing[1][44].t_rxd2[0][2] = 3295ns;
slave_timing[1][44].t_rxd2[2][0] = 1275ns;
slave_timing[1][44].t_rxd2[1][2] = 2898ns;
slave_timing[1][44].t_rxd2[2][1] = 1607ns;

slave_timing[1][45].info_corner          = 0;
slave_timing[1][45].info_temp__j__       = 25;
slave_timing[1][45].info_i__quite_rec__  = 0.000000000;
slave_timing[1][45].info_dtr__ib__       = 1;
slave_timing[1][45].info_i__offset_rec__ = 0.001000000;
slave_timing[1][45].info_i__max_slave__  = 0.021000000;
slave_timing[1][45].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][45].info_r__dsi_bus__    = 5.000;

slave_timing[1][45].t_rxd1[0][1] = 2125ns;
slave_timing[1][45].t_rxd1[1][0] = 1996ns;
slave_timing[1][45].t_rxd1[0][2] = 1570ns;
slave_timing[1][45].t_rxd1[2][0] = 2384ns;
slave_timing[1][45].t_rxd2[0][2] = 2596ns;
slave_timing[1][45].t_rxd2[2][0] = 1467ns;
slave_timing[1][45].t_rxd2[1][2] = 2273ns;
slave_timing[1][45].t_rxd2[2][1] = 1898ns;

slave_timing[1][46].info_corner          = 0;
slave_timing[1][46].info_temp__j__       = 25;
slave_timing[1][46].info_i__quite_rec__  = 0.000000000;
slave_timing[1][46].info_dtr__ib__       = 1;
slave_timing[1][46].info_i__offset_rec__ = -0.001000000;
slave_timing[1][46].info_i__max_slave__  = 0.027000000;
slave_timing[1][46].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][46].info_r__dsi_bus__    = 5.000;

slave_timing[1][46].t_rxd1[0][1] = 2123ns;
slave_timing[1][46].t_rxd1[1][0] = 1869ns;
slave_timing[1][46].t_rxd1[0][2] = 1577ns;
slave_timing[1][46].t_rxd1[2][0] = 2286ns;
slave_timing[1][46].t_rxd2[0][2] = 2282ns;
slave_timing[1][46].t_rxd2[2][0] = 1591ns;
slave_timing[1][46].t_rxd2[1][2] = 1847ns;
slave_timing[1][46].t_rxd2[2][1] = 2190ns;

slave_timing[1][47].info_corner          = 0;
slave_timing[1][47].info_temp__j__       = 25;
slave_timing[1][47].info_i__quite_rec__  = 0.000000000;
slave_timing[1][47].info_dtr__ib__       = 1;
slave_timing[1][47].info_i__offset_rec__ = 0.001000000;
slave_timing[1][47].info_i__max_slave__  = 0.027000000;
slave_timing[1][47].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][47].info_r__dsi_bus__    = 5.000;

slave_timing[1][47].t_rxd1[0][1] = 1872ns;
slave_timing[1][47].t_rxd1[1][0] = 2142ns;
slave_timing[1][47].t_rxd1[0][2] = 1444ns;
slave_timing[1][47].t_rxd1[2][0] = 2501ns;
slave_timing[1][47].t_rxd2[0][2] = 2118ns;
slave_timing[1][47].t_rxd2[2][0] = 1715ns;
slave_timing[1][47].t_rxd2[1][2] = 1644ns;
slave_timing[1][47].t_rxd2[2][1] = 2524ns;

slave_timing[1][48].info_corner          = 0;
slave_timing[1][48].info_temp__j__       = 25;
slave_timing[1][48].info_i__quite_rec__  = 0.040000000;
slave_timing[1][48].info_dtr__ib__       = -1;
slave_timing[1][48].info_i__offset_rec__ = -0.001000000;
slave_timing[1][48].info_i__max_slave__  = 0.021000000;
slave_timing[1][48].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][48].info_r__dsi_bus__    = 5.000;

slave_timing[1][48].t_rxd1[0][1] = 2039ns;
slave_timing[1][48].t_rxd1[1][0] = 1632ns;
slave_timing[1][48].t_rxd1[0][2] = 1443ns;
slave_timing[1][48].t_rxd1[2][0] = 2015ns;
slave_timing[1][48].t_rxd2[0][2] = 2337ns;
slave_timing[1][48].t_rxd2[2][0] = 1262ns;
slave_timing[1][48].t_rxd2[1][2] = 2058ns;
slave_timing[1][48].t_rxd2[2][1] = 1632ns;

slave_timing[1][49].info_corner          = 0;
slave_timing[1][49].info_temp__j__       = 25;
slave_timing[1][49].info_i__quite_rec__  = 0.040000000;
slave_timing[1][49].info_dtr__ib__       = -1;
slave_timing[1][49].info_i__offset_rec__ = 0.001000000;
slave_timing[1][49].info_i__max_slave__  = 0.021000000;
slave_timing[1][49].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][49].info_r__dsi_bus__    = 5.000;

slave_timing[1][49].t_rxd1[0][1] = 1723ns;
slave_timing[1][49].t_rxd1[1][0] = 1921ns;
slave_timing[1][49].t_rxd1[0][2] = 1304ns;
slave_timing[1][49].t_rxd1[2][0] = 2233ns;
slave_timing[1][49].t_rxd2[0][2] = 2085ns;
slave_timing[1][49].t_rxd2[2][0] = 1404ns;
slave_timing[1][49].t_rxd2[1][2] = 1736ns;
slave_timing[1][49].t_rxd2[2][1] = 1920ns;

slave_timing[1][50].info_corner          = 0;
slave_timing[1][50].info_temp__j__       = 25;
slave_timing[1][50].info_i__quite_rec__  = 0.040000000;
slave_timing[1][50].info_dtr__ib__       = -1;
slave_timing[1][50].info_i__offset_rec__ = -0.001000000;
slave_timing[1][50].info_i__max_slave__  = 0.027000000;
slave_timing[1][50].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][50].info_r__dsi_bus__    = 5.000;

slave_timing[1][50].t_rxd1[0][1] = 1796ns;
slave_timing[1][50].t_rxd1[1][0] = 1744ns;
slave_timing[1][50].t_rxd1[0][2] = 1339ns;
slave_timing[1][50].t_rxd1[2][0] = 2093ns;
slave_timing[1][50].t_rxd2[0][2] = 1917ns;
slave_timing[1][50].t_rxd2[2][0] = 1478ns;
slave_timing[1][50].t_rxd2[1][2] = 1490ns;
slave_timing[1][50].t_rxd2[2][1] = 2132ns;

slave_timing[1][51].info_corner          = 0;
slave_timing[1][51].info_temp__j__       = 25;
slave_timing[1][51].info_i__quite_rec__  = 0.040000000;
slave_timing[1][51].info_dtr__ib__       = -1;
slave_timing[1][51].info_i__offset_rec__ = 0.001000000;
slave_timing[1][51].info_i__max_slave__  = 0.027000000;
slave_timing[1][51].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][51].info_r__dsi_bus__    = 5.000;

slave_timing[1][51].t_rxd1[0][1] = 1601ns;
slave_timing[1][51].t_rxd1[1][0] = 1957ns;
slave_timing[1][51].t_rxd1[0][2] = 1223ns;
slave_timing[1][51].t_rxd1[2][0] = 2264ns;
slave_timing[1][51].t_rxd2[0][2] = 1796ns;
slave_timing[1][51].t_rxd2[2][0] = 1569ns;
slave_timing[1][51].t_rxd2[1][2] = 1297ns;
slave_timing[1][51].t_rxd2[2][1] = 2636ns;

slave_timing[1][52].info_corner          = 0;
slave_timing[1][52].info_temp__j__       = 25;
slave_timing[1][52].info_i__quite_rec__  = 0.040000000;
slave_timing[1][52].info_dtr__ib__       = 1;
slave_timing[1][52].info_i__offset_rec__ = -0.001000000;
slave_timing[1][52].info_i__max_slave__  = 0.021000000;
slave_timing[1][52].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][52].info_r__dsi_bus__    = 5.000;

slave_timing[1][52].t_rxd1[0][1] = 2309ns;
slave_timing[1][52].t_rxd1[1][0] = 1496ns;
slave_timing[1][52].t_rxd1[0][2] = 1521ns;
slave_timing[1][52].t_rxd1[2][0] = 1926ns;
slave_timing[1][52].t_rxd2[0][2] = 2848ns;
slave_timing[1][52].t_rxd2[2][0] = 1123ns;
slave_timing[1][52].t_rxd2[1][2] = 2615ns;
slave_timing[1][52].t_rxd2[2][1] = 1410ns;

slave_timing[1][53].info_corner          = 0;
slave_timing[1][53].info_temp__j__       = 25;
slave_timing[1][53].info_i__quite_rec__  = 0.040000000;
slave_timing[1][53].info_dtr__ib__       = 1;
slave_timing[1][53].info_i__offset_rec__ = 0.001000000;
slave_timing[1][53].info_i__max_slave__  = 0.021000000;
slave_timing[1][53].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][53].info_r__dsi_bus__    = 5.000;

slave_timing[1][53].t_rxd1[0][1] = 1900ns;
slave_timing[1][53].t_rxd1[1][0] = 1766ns;
slave_timing[1][53].t_rxd1[0][2] = 1384ns;
slave_timing[1][53].t_rxd1[2][0] = 2110ns;
slave_timing[1][53].t_rxd2[0][2] = 2315ns;
slave_timing[1][53].t_rxd2[2][0] = 1285ns;
slave_timing[1][53].t_rxd2[1][2] = 2034ns;
slave_timing[1][53].t_rxd2[2][1] = 1678ns;

slave_timing[1][54].info_corner          = 0;
slave_timing[1][54].info_temp__j__       = 25;
slave_timing[1][54].info_i__quite_rec__  = 0.040000000;
slave_timing[1][54].info_dtr__ib__       = 1;
slave_timing[1][54].info_i__offset_rec__ = -0.001000000;
slave_timing[1][54].info_i__max_slave__  = 0.027000000;
slave_timing[1][54].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][54].info_r__dsi_bus__    = 5.000;

slave_timing[1][54].t_rxd1[0][1] = 1919ns;
slave_timing[1][54].t_rxd1[1][0] = 1651ns;
slave_timing[1][54].t_rxd1[0][2] = 1393ns;
slave_timing[1][54].t_rxd1[2][0] = 2026ns;
slave_timing[1][54].t_rxd2[0][2] = 2033ns;
slave_timing[1][54].t_rxd2[2][0] = 1399ns;
slave_timing[1][54].t_rxd2[1][2] = 1665ns;
slave_timing[1][54].t_rxd2[2][1] = 1916ns;

slave_timing[1][55].info_corner          = 0;
slave_timing[1][55].info_temp__j__       = 25;
slave_timing[1][55].info_i__quite_rec__  = 0.040000000;
slave_timing[1][55].info_dtr__ib__       = 1;
slave_timing[1][55].info_i__offset_rec__ = 0.001000000;
slave_timing[1][55].info_i__max_slave__  = 0.027000000;
slave_timing[1][55].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][55].info_r__dsi_bus__    = 5.000;

slave_timing[1][55].t_rxd1[0][1] = 1688ns;
slave_timing[1][55].t_rxd1[1][0] = 1872ns;
slave_timing[1][55].t_rxd1[0][2] = 1283ns;
slave_timing[1][55].t_rxd1[2][0] = 2192ns;
slave_timing[1][55].t_rxd2[0][2] = 1896ns;
slave_timing[1][55].t_rxd2[2][0] = 1503ns;
slave_timing[1][55].t_rxd2[1][2] = 1455ns;
slave_timing[1][55].t_rxd2[2][1] = 2224ns;

slave_timing[1][56].info_corner          = 0;
slave_timing[1][56].info_temp__j__       = 25;
slave_timing[1][56].info_i__quite_rec__  = 0.040000000;
slave_timing[1][56].info_dtr__ib__       = -1;
slave_timing[1][56].info_i__offset_rec__ = -0.001000000;
slave_timing[1][56].info_i__max_slave__  = 0.021000000;
slave_timing[1][56].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][56].info_r__dsi_bus__    = 5.000;

slave_timing[1][56].t_rxd1[0][1] = 2289ns;
slave_timing[1][56].t_rxd1[1][0] = 1840ns;
slave_timing[1][56].t_rxd1[0][2] = 1634ns;
slave_timing[1][56].t_rxd1[2][0] = 2266ns;
slave_timing[1][56].t_rxd2[0][2] = 2628ns;
slave_timing[1][56].t_rxd2[2][0] = 1438ns;
slave_timing[1][56].t_rxd2[1][2] = 2310ns;
slave_timing[1][56].t_rxd2[2][1] = 1843ns;

slave_timing[1][57].info_corner          = 0;
slave_timing[1][57].info_temp__j__       = 25;
slave_timing[1][57].info_i__quite_rec__  = 0.040000000;
slave_timing[1][57].info_dtr__ib__       = -1;
slave_timing[1][57].info_i__offset_rec__ = 0.001000000;
slave_timing[1][57].info_i__max_slave__  = 0.021000000;
slave_timing[1][57].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][57].info_r__dsi_bus__    = 5.000;

slave_timing[1][57].t_rxd1[0][1] = 1943ns;
slave_timing[1][57].t_rxd1[1][0] = 2157ns;
slave_timing[1][57].t_rxd1[0][2] = 1485ns;
slave_timing[1][57].t_rxd1[2][0] = 2516ns;
slave_timing[1][57].t_rxd2[0][2] = 2345ns;
slave_timing[1][57].t_rxd2[2][0] = 1594ns;
slave_timing[1][57].t_rxd2[1][2] = 1957ns;
slave_timing[1][57].t_rxd2[2][1] = 2160ns;

slave_timing[1][58].info_corner          = 0;
slave_timing[1][58].info_temp__j__       = 25;
slave_timing[1][58].info_i__quite_rec__  = 0.040000000;
slave_timing[1][58].info_dtr__ib__       = -1;
slave_timing[1][58].info_i__offset_rec__ = -0.001000000;
slave_timing[1][58].info_i__max_slave__  = 0.027000000;
slave_timing[1][58].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][58].info_r__dsi_bus__    = 5.000;

slave_timing[1][58].t_rxd1[0][1] = 2024ns;
slave_timing[1][58].t_rxd1[1][0] = 1962ns;
slave_timing[1][58].t_rxd1[0][2] = 1521ns;
slave_timing[1][58].t_rxd1[2][0] = 2356ns;
slave_timing[1][58].t_rxd2[0][2] = 2156ns;
slave_timing[1][58].t_rxd2[2][0] = 1675ns;
slave_timing[1][58].t_rxd2[1][2] = 1684ns;
slave_timing[1][58].t_rxd2[2][1] = 2402ns;

slave_timing[1][59].info_corner          = 0;
slave_timing[1][59].info_temp__j__       = 25;
slave_timing[1][59].info_i__quite_rec__  = 0.040000000;
slave_timing[1][59].info_dtr__ib__       = -1;
slave_timing[1][59].info_i__offset_rec__ = 0.001000000;
slave_timing[1][59].info_i__max_slave__  = 0.027000000;
slave_timing[1][59].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][59].info_r__dsi_bus__    = 5.000;

slave_timing[1][59].t_rxd1[0][1] = 1808ns;
slave_timing[1][59].t_rxd1[1][0] = 2202ns;
slave_timing[1][59].t_rxd1[0][2] = 1396ns;
slave_timing[1][59].t_rxd1[2][0] = 2550ns;
slave_timing[1][59].t_rxd2[0][2] = 2022ns;
slave_timing[1][59].t_rxd2[2][0] = 1773ns;
slave_timing[1][59].t_rxd2[1][2] = 1475ns;
slave_timing[1][59].t_rxd2[2][1] = 2973ns;

slave_timing[1][60].info_corner          = 0;
slave_timing[1][60].info_temp__j__       = 25;
slave_timing[1][60].info_i__quite_rec__  = 0.040000000;
slave_timing[1][60].info_dtr__ib__       = 1;
slave_timing[1][60].info_i__offset_rec__ = -0.001000000;
slave_timing[1][60].info_i__max_slave__  = 0.021000000;
slave_timing[1][60].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][60].info_r__dsi_bus__    = 5.000;

slave_timing[1][60].t_rxd1[0][1] = 2591ns;
slave_timing[1][60].t_rxd1[1][0] = 1693ns;
slave_timing[1][60].t_rxd1[0][2] = 1722ns;
slave_timing[1][60].t_rxd1[2][0] = 2167ns;
slave_timing[1][60].t_rxd2[0][2] = 3201ns;
slave_timing[1][60].t_rxd2[2][0] = 1291ns;
slave_timing[1][60].t_rxd2[1][2] = 2947ns;
slave_timing[1][60].t_rxd2[2][1] = 1598ns;

slave_timing[1][61].info_corner          = 0;
slave_timing[1][61].info_temp__j__       = 25;
slave_timing[1][61].info_i__quite_rec__  = 0.040000000;
slave_timing[1][61].info_dtr__ib__       = 1;
slave_timing[1][61].info_i__offset_rec__ = 0.001000000;
slave_timing[1][61].info_i__max_slave__  = 0.021000000;
slave_timing[1][61].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][61].info_r__dsi_bus__    = 5.000;

slave_timing[1][61].t_rxd1[0][1] = 2136ns;
slave_timing[1][61].t_rxd1[1][0] = 1986ns;
slave_timing[1][61].t_rxd1[0][2] = 1574ns;
slave_timing[1][61].t_rxd1[2][0] = 2377ns;
slave_timing[1][61].t_rxd2[0][2] = 2606ns;
slave_timing[1][61].t_rxd2[2][0] = 1465ns;
slave_timing[1][61].t_rxd2[1][2] = 2286ns;
slave_timing[1][61].t_rxd2[2][1] = 1891ns;

slave_timing[1][62].info_corner          = 0;
slave_timing[1][62].info_temp__j__       = 25;
slave_timing[1][62].info_i__quite_rec__  = 0.040000000;
slave_timing[1][62].info_dtr__ib__       = 1;
slave_timing[1][62].info_i__offset_rec__ = -0.001000000;
slave_timing[1][62].info_i__max_slave__  = 0.027000000;
slave_timing[1][62].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][62].info_r__dsi_bus__    = 5.000;

slave_timing[1][62].t_rxd1[0][1] = 2159ns;
slave_timing[1][62].t_rxd1[1][0] = 1860ns;
slave_timing[1][62].t_rxd1[0][2] = 1582ns;
slave_timing[1][62].t_rxd1[2][0] = 2280ns;
slave_timing[1][62].t_rxd2[0][2] = 2286ns;
slave_timing[1][62].t_rxd2[2][0] = 1588ns;
slave_timing[1][62].t_rxd2[1][2] = 1878ns;
slave_timing[1][62].t_rxd2[2][1] = 2154ns;

slave_timing[1][63].info_corner          = 0;
slave_timing[1][63].info_temp__j__       = 25;
slave_timing[1][63].info_i__quite_rec__  = 0.040000000;
slave_timing[1][63].info_dtr__ib__       = 1;
slave_timing[1][63].info_i__offset_rec__ = 0.001000000;
slave_timing[1][63].info_i__max_slave__  = 0.027000000;
slave_timing[1][63].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][63].info_r__dsi_bus__    = 5.000;

slave_timing[1][63].t_rxd1[0][1] = 1906ns;
slave_timing[1][63].t_rxd1[1][0] = 2107ns;
slave_timing[1][63].t_rxd1[0][2] = 1462ns;
slave_timing[1][63].t_rxd1[2][0] = 2469ns;
slave_timing[1][63].t_rxd2[0][2] = 2134ns;
slave_timing[1][63].t_rxd2[2][0] = 1703ns;
slave_timing[1][63].t_rxd2[1][2] = 1650ns;
slave_timing[1][63].t_rxd2[2][1] = 2508ns;

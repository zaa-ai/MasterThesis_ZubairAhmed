
slave_timing[0][32+0].info_corner          = 2;
slave_timing[0][32+0].info_temp__j__       = 125;
slave_timing[0][32+0].info_i__quite_rec__  = 0.006000000;
slave_timing[0][32+0].info_dtr__ib__       = -1;
slave_timing[0][32+0].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+0].info_i__max_slave__  = 0.023000000;
slave_timing[0][32+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][32+0].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+0].t_rxd1[0][1] = 1109ns;
slave_timing[0][32+0].t_rxd1[1][0] = 1136ns;
slave_timing[0][32+0].t_rxd1[0][2] = 823ns;
slave_timing[0][32+0].t_rxd1[2][0] = 1398ns;
slave_timing[0][32+0].t_rxd2[0][2] = 1355ns;
slave_timing[0][32+0].t_rxd2[2][0] = 836ns;
slave_timing[0][32+0].t_rxd2[1][2] = 1095ns;
slave_timing[0][32+0].t_rxd2[2][1] = 1116ns;

slave_timing[0][32+1].info_corner          = 2;
slave_timing[0][32+1].info_temp__j__       = 125;
slave_timing[0][32+1].info_i__quite_rec__  = 0.006000000;
slave_timing[0][32+1].info_dtr__ib__       = -1;
slave_timing[0][32+1].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+1].info_i__max_slave__  = 0.025000000;
slave_timing[0][32+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][32+1].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+1].t_rxd1[0][1] = 1062ns;
slave_timing[0][32+1].t_rxd1[1][0] = 1168ns;
slave_timing[0][32+1].t_rxd1[0][2] = 801ns;
slave_timing[0][32+1].t_rxd1[2][0] = 1428ns;
slave_timing[0][32+1].t_rxd2[0][2] = 1258ns;
slave_timing[0][32+1].t_rxd2[2][0] = 888ns;
slave_timing[0][32+1].t_rxd2[1][2] = 971ns;
slave_timing[0][32+1].t_rxd2[2][1] = 1243ns;

slave_timing[0][32+2].info_corner          = 2;
slave_timing[0][32+2].info_temp__j__       = 125;
slave_timing[0][32+2].info_i__quite_rec__  = 0.006000000;
slave_timing[0][32+2].info_dtr__ib__       = 1;
slave_timing[0][32+2].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+2].info_i__max_slave__  = 0.023000000;
slave_timing[0][32+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][32+2].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+2].t_rxd1[0][1] = 1128ns;
slave_timing[0][32+2].t_rxd1[1][0] = 1101ns;
slave_timing[0][32+2].t_rxd1[0][2] = 828ns;
slave_timing[0][32+2].t_rxd1[2][0] = 1363ns;
slave_timing[0][32+2].t_rxd2[0][2] = 1436ns;
slave_timing[0][32+2].t_rxd2[2][0] = 788ns;
slave_timing[0][32+2].t_rxd2[1][2] = 1197ns;
slave_timing[0][32+2].t_rxd2[2][1] = 1019ns;

slave_timing[0][32+3].info_corner          = 2;
slave_timing[0][32+3].info_temp__j__       = 125;
slave_timing[0][32+3].info_i__quite_rec__  = 0.006000000;
slave_timing[0][32+3].info_dtr__ib__       = 1;
slave_timing[0][32+3].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+3].info_i__max_slave__  = 0.025000000;
slave_timing[0][32+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][32+3].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+3].t_rxd1[0][1] = 1079ns;
slave_timing[0][32+3].t_rxd1[1][0] = 1136ns;
slave_timing[0][32+3].t_rxd1[0][2] = 803ns;
slave_timing[0][32+3].t_rxd1[2][0] = 1391ns;
slave_timing[0][32+3].t_rxd2[0][2] = 1312ns;
slave_timing[0][32+3].t_rxd2[2][0] = 844ns;
slave_timing[0][32+3].t_rxd2[1][2] = 1055ns;
slave_timing[0][32+3].t_rxd2[2][1] = 1135ns;

slave_timing[0][32+4].info_corner          = 2;
slave_timing[0][32+4].info_temp__j__       = 125;
slave_timing[0][32+4].info_i__quite_rec__  = 0.006000000;
slave_timing[0][32+4].info_dtr__ib__       = -1;
slave_timing[0][32+4].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+4].info_i__max_slave__  = 0.023000000;
slave_timing[0][32+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][32+4].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+4].t_rxd1[0][1] = 1279ns;
slave_timing[0][32+4].t_rxd1[1][0] = 1269ns;
slave_timing[0][32+4].t_rxd1[0][2] = 946ns;
slave_timing[0][32+4].t_rxd1[2][0] = 1519ns;
slave_timing[0][32+4].t_rxd2[0][2] = 1407ns;
slave_timing[0][32+4].t_rxd2[2][0] = 872ns;
slave_timing[0][32+4].t_rxd2[1][2] = 1117ns;
slave_timing[0][32+4].t_rxd2[2][1] = 1139ns;

slave_timing[0][32+5].info_corner          = 2;
slave_timing[0][32+5].info_temp__j__       = 125;
slave_timing[0][32+5].info_i__quite_rec__  = 0.006000000;
slave_timing[0][32+5].info_dtr__ib__       = -1;
slave_timing[0][32+5].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+5].info_i__max_slave__  = 0.025000000;
slave_timing[0][32+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][32+5].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+5].t_rxd1[0][1] = 1223ns;
slave_timing[0][32+5].t_rxd1[1][0] = 1303ns;
slave_timing[0][32+5].t_rxd1[0][2] = 919ns;
slave_timing[0][32+5].t_rxd1[2][0] = 1547ns;
slave_timing[0][32+5].t_rxd2[0][2] = 1311ns;
slave_timing[0][32+5].t_rxd2[2][0] = 924ns;
slave_timing[0][32+5].t_rxd2[1][2] = 1000ns;
slave_timing[0][32+5].t_rxd2[2][1] = 1260ns;

slave_timing[0][32+6].info_corner          = 2;
slave_timing[0][32+6].info_temp__j__       = 125;
slave_timing[0][32+6].info_i__quite_rec__  = 0.006000000;
slave_timing[0][32+6].info_dtr__ib__       = 1;
slave_timing[0][32+6].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+6].info_i__max_slave__  = 0.023000000;
slave_timing[0][32+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][32+6].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+6].t_rxd1[0][1] = 1304ns;
slave_timing[0][32+6].t_rxd1[1][0] = 1231ns;
slave_timing[0][32+6].t_rxd1[0][2] = 954ns;
slave_timing[0][32+6].t_rxd1[2][0] = 1485ns;
slave_timing[0][32+6].t_rxd2[0][2] = 1485ns;
slave_timing[0][32+6].t_rxd2[2][0] = 824ns;
slave_timing[0][32+6].t_rxd2[1][2] = 1213ns;
slave_timing[0][32+6].t_rxd2[2][1] = 1043ns;

slave_timing[0][32+7].info_corner          = 2;
slave_timing[0][32+7].info_temp__j__       = 125;
slave_timing[0][32+7].info_i__quite_rec__  = 0.006000000;
slave_timing[0][32+7].info_dtr__ib__       = 1;
slave_timing[0][32+7].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+7].info_i__max_slave__  = 0.025000000;
slave_timing[0][32+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][32+7].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+7].t_rxd1[0][1] = 1243ns;
slave_timing[0][32+7].t_rxd1[1][0] = 1267ns;
slave_timing[0][32+7].t_rxd1[0][2] = 926ns;
slave_timing[0][32+7].t_rxd1[2][0] = 1509ns;
slave_timing[0][32+7].t_rxd2[0][2] = 1362ns;
slave_timing[0][32+7].t_rxd2[2][0] = 876ns;
slave_timing[0][32+7].t_rxd2[1][2] = 1076ns;
slave_timing[0][32+7].t_rxd2[2][1] = 1141ns;

slave_timing[0][32+8].info_corner          = 2;
slave_timing[0][32+8].info_temp__j__       = 125;
slave_timing[0][32+8].info_i__quite_rec__  = 0.003000000;
slave_timing[0][32+8].info_dtr__ib__       = -1;
slave_timing[0][32+8].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+8].info_i__max_slave__  = 0.023000000;
slave_timing[0][32+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][32+8].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+8].t_rxd1[0][1] = 1093ns;
slave_timing[0][32+8].t_rxd1[1][0] = 1113ns;
slave_timing[0][32+8].t_rxd1[0][2] = 814ns;
slave_timing[0][32+8].t_rxd1[2][0] = 1369ns;
slave_timing[0][32+8].t_rxd2[0][2] = 1339ns;
slave_timing[0][32+8].t_rxd2[2][0] = 827ns;
slave_timing[0][32+8].t_rxd2[1][2] = 1093ns;
slave_timing[0][32+8].t_rxd2[2][1] = 1097ns;

slave_timing[0][32+9].info_corner          = 2;
slave_timing[0][32+9].info_temp__j__       = 125;
slave_timing[0][32+9].info_i__quite_rec__  = 0.003000000;
slave_timing[0][32+9].info_dtr__ib__       = -1;
slave_timing[0][32+9].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+9].info_i__max_slave__  = 0.025000000;
slave_timing[0][32+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][32+9].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+9].t_rxd1[0][1] = 1046ns;
slave_timing[0][32+9].t_rxd1[1][0] = 1144ns;
slave_timing[0][32+9].t_rxd1[0][2] = 789ns;
slave_timing[0][32+9].t_rxd1[2][0] = 1397ns;
slave_timing[0][32+9].t_rxd2[0][2] = 1241ns;
slave_timing[0][32+9].t_rxd2[2][0] = 877ns;
slave_timing[0][32+9].t_rxd2[1][2] = 972ns;
slave_timing[0][32+9].t_rxd2[2][1] = 1221ns;

slave_timing[0][32+10].info_corner          = 2;
slave_timing[0][32+10].info_temp__j__       = 125;
slave_timing[0][32+10].info_i__quite_rec__  = 0.003000000;
slave_timing[0][32+10].info_dtr__ib__       = 1;
slave_timing[0][32+10].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+10].info_i__max_slave__  = 0.023000000;
slave_timing[0][32+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][32+10].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+10].t_rxd1[0][1] = 1104ns;
slave_timing[0][32+10].t_rxd1[1][0] = 1067ns;
slave_timing[0][32+10].t_rxd1[0][2] = 813ns;
slave_timing[0][32+10].t_rxd1[2][0] = 1317ns;
slave_timing[0][32+10].t_rxd2[0][2] = 1413ns;
slave_timing[0][32+10].t_rxd2[2][0] = 777ns;
slave_timing[0][32+10].t_rxd2[1][2] = 1190ns;
slave_timing[0][32+10].t_rxd2[2][1] = 1002ns;

slave_timing[0][32+11].info_corner          = 2;
slave_timing[0][32+11].info_temp__j__       = 125;
slave_timing[0][32+11].info_i__quite_rec__  = 0.003000000;
slave_timing[0][32+11].info_dtr__ib__       = 1;
slave_timing[0][32+11].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+11].info_i__max_slave__  = 0.025000000;
slave_timing[0][32+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][32+11].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+11].t_rxd1[0][1] = 1055ns;
slave_timing[0][32+11].t_rxd1[1][0] = 1098ns;
slave_timing[0][32+11].t_rxd1[0][2] = 790ns;
slave_timing[0][32+11].t_rxd1[2][0] = 1344ns;
slave_timing[0][32+11].t_rxd2[0][2] = 1291ns;
slave_timing[0][32+11].t_rxd2[2][0] = 833ns;
slave_timing[0][32+11].t_rxd2[1][2] = 1049ns;
slave_timing[0][32+11].t_rxd2[2][1] = 1117ns;

slave_timing[0][32+12].info_corner          = 2;
slave_timing[0][32+12].info_temp__j__       = 125;
slave_timing[0][32+12].info_i__quite_rec__  = 0.003000000;
slave_timing[0][32+12].info_dtr__ib__       = -1;
slave_timing[0][32+12].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+12].info_i__max_slave__  = 0.023000000;
slave_timing[0][32+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][32+12].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+12].t_rxd1[0][1] = 1277ns;
slave_timing[0][32+12].t_rxd1[1][0] = 1248ns;
slave_timing[0][32+12].t_rxd1[0][2] = 945ns;
slave_timing[0][32+12].t_rxd1[2][0] = 1489ns;
slave_timing[0][32+12].t_rxd2[0][2] = 1389ns;
slave_timing[0][32+12].t_rxd2[2][0] = 861ns;
slave_timing[0][32+12].t_rxd2[1][2] = 1113ns;
slave_timing[0][32+12].t_rxd2[2][1] = 1118ns;

slave_timing[0][32+13].info_corner          = 2;
slave_timing[0][32+13].info_temp__j__       = 125;
slave_timing[0][32+13].info_i__quite_rec__  = 0.003000000;
slave_timing[0][32+13].info_dtr__ib__       = -1;
slave_timing[0][32+13].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+13].info_i__max_slave__  = 0.025000000;
slave_timing[0][32+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][32+13].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+13].t_rxd1[0][1] = 1221ns;
slave_timing[0][32+13].t_rxd1[1][0] = 1280ns;
slave_timing[0][32+13].t_rxd1[0][2] = 917ns;
slave_timing[0][32+13].t_rxd1[2][0] = 1516ns;
slave_timing[0][32+13].t_rxd2[0][2] = 1293ns;
slave_timing[0][32+13].t_rxd2[2][0] = 912ns;
slave_timing[0][32+13].t_rxd2[1][2] = 997ns;
slave_timing[0][32+13].t_rxd2[2][1] = 1234ns;

slave_timing[0][32+14].info_corner          = 2;
slave_timing[0][32+14].info_temp__j__       = 125;
slave_timing[0][32+14].info_i__quite_rec__  = 0.003000000;
slave_timing[0][32+14].info_dtr__ib__       = 1;
slave_timing[0][32+14].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+14].info_i__max_slave__  = 0.023000000;
slave_timing[0][32+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][32+14].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+14].t_rxd1[0][1] = 1296ns;
slave_timing[0][32+14].t_rxd1[1][0] = 1195ns;
slave_timing[0][32+14].t_rxd1[0][2] = 948ns;
slave_timing[0][32+14].t_rxd1[2][0] = 1434ns;
slave_timing[0][32+14].t_rxd2[0][2] = 1460ns;
slave_timing[0][32+14].t_rxd2[2][0] = 811ns;
slave_timing[0][32+14].t_rxd2[1][2] = 1201ns;
slave_timing[0][32+14].t_rxd2[2][1] = 1024ns;

slave_timing[0][32+15].info_corner          = 2;
slave_timing[0][32+15].info_temp__j__       = 125;
slave_timing[0][32+15].info_i__quite_rec__  = 0.003000000;
slave_timing[0][32+15].info_dtr__ib__       = 1;
slave_timing[0][32+15].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+15].info_i__max_slave__  = 0.025000000;
slave_timing[0][32+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][32+15].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+15].t_rxd1[0][1] = 1236ns;
slave_timing[0][32+15].t_rxd1[1][0] = 1227ns;
slave_timing[0][32+15].t_rxd1[0][2] = 920ns;
slave_timing[0][32+15].t_rxd1[2][0] = 1461ns;
slave_timing[0][32+15].t_rxd2[0][2] = 1341ns;
slave_timing[0][32+15].t_rxd2[2][0] = 868ns;
slave_timing[0][32+15].t_rxd2[1][2] = 1069ns;
slave_timing[0][32+15].t_rxd2[2][1] = 1137ns;

slave_timing[0][32+16].info_corner          = 2;
slave_timing[0][32+16].info_temp__j__       = 125;
slave_timing[0][32+16].info_i__quite_rec__  = 0.000000000;
slave_timing[0][32+16].info_dtr__ib__       = -1;
slave_timing[0][32+16].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+16].info_i__max_slave__  = 0.023000000;
slave_timing[0][32+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][32+16].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+16].t_rxd1[0][1] = 1067ns;
slave_timing[0][32+16].t_rxd1[1][0] = 1081ns;
slave_timing[0][32+16].t_rxd1[0][2] = 796ns;
slave_timing[0][32+16].t_rxd1[2][0] = 1321ns;
slave_timing[0][32+16].t_rxd2[0][2] = 1310ns;
slave_timing[0][32+16].t_rxd2[2][0] = 812ns;
slave_timing[0][32+16].t_rxd2[1][2] = 1081ns;
slave_timing[0][32+16].t_rxd2[2][1] = 1077ns;

slave_timing[0][32+17].info_corner          = 2;
slave_timing[0][32+17].info_temp__j__       = 125;
slave_timing[0][32+17].info_i__quite_rec__  = 0.000000000;
slave_timing[0][32+17].info_dtr__ib__       = -1;
slave_timing[0][32+17].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+17].info_i__max_slave__  = 0.025000000;
slave_timing[0][32+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][32+17].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+17].t_rxd1[0][1] = 1021ns;
slave_timing[0][32+17].t_rxd1[1][0] = 1110ns;
slave_timing[0][32+17].t_rxd1[0][2] = 772ns;
slave_timing[0][32+17].t_rxd1[2][0] = 1347ns;
slave_timing[0][32+17].t_rxd2[0][2] = 1215ns;
slave_timing[0][32+17].t_rxd2[2][0] = 864ns;
slave_timing[0][32+17].t_rxd2[1][2] = 963ns;
slave_timing[0][32+17].t_rxd2[2][1] = 1196ns;

slave_timing[0][32+18].info_corner          = 2;
slave_timing[0][32+18].info_temp__j__       = 125;
slave_timing[0][32+18].info_i__quite_rec__  = 0.000000000;
slave_timing[0][32+18].info_dtr__ib__       = 1;
slave_timing[0][32+18].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+18].info_i__max_slave__  = 0.023000000;
slave_timing[0][32+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][32+18].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+18].t_rxd1[0][1] = 1078ns;
slave_timing[0][32+18].t_rxd1[1][0] = 1040ns;
slave_timing[0][32+18].t_rxd1[0][2] = 796ns;
slave_timing[0][32+18].t_rxd1[2][0] = 1274ns;
slave_timing[0][32+18].t_rxd2[0][2] = 1374ns;
slave_timing[0][32+18].t_rxd2[2][0] = 761ns;
slave_timing[0][32+18].t_rxd2[1][2] = 1166ns;
slave_timing[0][32+18].t_rxd2[2][1] = 973ns;

slave_timing[0][32+19].info_corner          = 2;
slave_timing[0][32+19].info_temp__j__       = 125;
slave_timing[0][32+19].info_i__quite_rec__  = 0.000000000;
slave_timing[0][32+19].info_dtr__ib__       = 1;
slave_timing[0][32+19].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+19].info_i__max_slave__  = 0.025000000;
slave_timing[0][32+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][32+19].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+19].t_rxd1[0][1] = 1031ns;
slave_timing[0][32+19].t_rxd1[1][0] = 1067ns;
slave_timing[0][32+19].t_rxd1[0][2] = 774ns;
slave_timing[0][32+19].t_rxd1[2][0] = 1300ns;
slave_timing[0][32+19].t_rxd2[0][2] = 1256ns;
slave_timing[0][32+19].t_rxd2[2][0] = 817ns;
slave_timing[0][32+19].t_rxd2[1][2] = 1031ns;
slave_timing[0][32+19].t_rxd2[2][1] = 1087ns;

slave_timing[0][32+20].info_corner          = 2;
slave_timing[0][32+20].info_temp__j__       = 125;
slave_timing[0][32+20].info_i__quite_rec__  = 0.000000000;
slave_timing[0][32+20].info_dtr__ib__       = -1;
slave_timing[0][32+20].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+20].info_i__max_slave__  = 0.023000000;
slave_timing[0][32+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][32+20].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+20].t_rxd1[0][1] = 1270ns;
slave_timing[0][32+20].t_rxd1[1][0] = 1206ns;
slave_timing[0][32+20].t_rxd1[0][2] = 940ns;
slave_timing[0][32+20].t_rxd1[2][0] = 1435ns;
slave_timing[0][32+20].t_rxd2[0][2] = 1356ns;
slave_timing[0][32+20].t_rxd2[2][0] = 849ns;
slave_timing[0][32+20].t_rxd2[1][2] = 1099ns;
slave_timing[0][32+20].t_rxd2[2][1] = 1083ns;

slave_timing[0][32+21].info_corner          = 2;
slave_timing[0][32+21].info_temp__j__       = 125;
slave_timing[0][32+21].info_i__quite_rec__  = 0.000000000;
slave_timing[0][32+21].info_dtr__ib__       = -1;
slave_timing[0][32+21].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+21].info_i__max_slave__  = 0.025000000;
slave_timing[0][32+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][32+21].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+21].t_rxd1[0][1] = 1214ns;
slave_timing[0][32+21].t_rxd1[1][0] = 1235ns;
slave_timing[0][32+21].t_rxd1[0][2] = 912ns;
slave_timing[0][32+21].t_rxd1[2][0] = 1459ns;
slave_timing[0][32+21].t_rxd2[0][2] = 1266ns;
slave_timing[0][32+21].t_rxd2[2][0] = 898ns;
slave_timing[0][32+21].t_rxd2[1][2] = 983ns;
slave_timing[0][32+21].t_rxd2[2][1] = 1207ns;

slave_timing[0][32+22].info_corner          = 2;
slave_timing[0][32+22].info_temp__j__       = 125;
slave_timing[0][32+22].info_i__quite_rec__  = 0.000000000;
slave_timing[0][32+22].info_dtr__ib__       = 1;
slave_timing[0][32+22].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+22].info_i__max_slave__  = 0.023000000;
slave_timing[0][32+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][32+22].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+22].t_rxd1[0][1] = 1291ns;
slave_timing[0][32+22].t_rxd1[1][0] = 1165ns;
slave_timing[0][32+22].t_rxd1[0][2] = 943ns;
slave_timing[0][32+22].t_rxd1[2][0] = 1386ns;
slave_timing[0][32+22].t_rxd2[0][2] = 1414ns;
slave_timing[0][32+22].t_rxd2[2][0] = 794ns;
slave_timing[0][32+22].t_rxd2[1][2] = 1181ns;
slave_timing[0][32+22].t_rxd2[2][1] = 985ns;

slave_timing[0][32+23].info_corner          = 2;
slave_timing[0][32+23].info_temp__j__       = 125;
slave_timing[0][32+23].info_i__quite_rec__  = 0.000000000;
slave_timing[0][32+23].info_dtr__ib__       = 1;
slave_timing[0][32+23].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+23].info_i__max_slave__  = 0.025000000;
slave_timing[0][32+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][32+23].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+23].t_rxd1[0][1] = 1231ns;
slave_timing[0][32+23].t_rxd1[1][0] = 1194ns;
slave_timing[0][32+23].t_rxd1[0][2] = 915ns;
slave_timing[0][32+23].t_rxd1[2][0] = 1412ns;
slave_timing[0][32+23].t_rxd2[0][2] = 1301ns;
slave_timing[0][32+23].t_rxd2[2][0] = 849ns;
slave_timing[0][32+23].t_rxd2[1][2] = 1050ns;
slave_timing[0][32+23].t_rxd2[2][1] = 1093ns;

slave_timing[0][32+24].info_corner          = 2;
slave_timing[0][32+24].info_temp__j__       = 125;
slave_timing[0][32+24].info_i__quite_rec__  = 0.040000000;
slave_timing[0][32+24].info_dtr__ib__       = -1;
slave_timing[0][32+24].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+24].info_i__max_slave__  = 0.023000000;
slave_timing[0][32+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][32+24].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+24].t_rxd1[0][1] = 1104ns;
slave_timing[0][32+24].t_rxd1[1][0] = 1136ns;
slave_timing[0][32+24].t_rxd1[0][2] = 833ns;
slave_timing[0][32+24].t_rxd1[2][0] = 1422ns;
slave_timing[0][32+24].t_rxd2[0][2] = 1525ns;
slave_timing[0][32+24].t_rxd2[2][0] = 980ns;
slave_timing[0][32+24].t_rxd2[1][2] = 1282ns;
slave_timing[0][32+24].t_rxd2[2][1] = 1310ns;

slave_timing[0][32+25].info_corner          = 2;
slave_timing[0][32+25].info_temp__j__       = 125;
slave_timing[0][32+25].info_i__quite_rec__  = 0.040000000;
slave_timing[0][32+25].info_dtr__ib__       = -1;
slave_timing[0][32+25].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+25].info_i__max_slave__  = 0.025000000;
slave_timing[0][32+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][32+25].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+25].t_rxd1[0][1] = 1058ns;
slave_timing[0][32+25].t_rxd1[1][0] = 1169ns;
slave_timing[0][32+25].t_rxd1[0][2] = 808ns;
slave_timing[0][32+25].t_rxd1[2][0] = 1458ns;
slave_timing[0][32+25].t_rxd2[0][2] = 1422ns;
slave_timing[0][32+25].t_rxd2[2][0] = 1033ns;
slave_timing[0][32+25].t_rxd2[1][2] = 1154ns;
slave_timing[0][32+25].t_rxd2[2][1] = 1441ns;

slave_timing[0][32+26].info_corner          = 2;
slave_timing[0][32+26].info_temp__j__       = 125;
slave_timing[0][32+26].info_i__quite_rec__  = 0.040000000;
slave_timing[0][32+26].info_dtr__ib__       = 1;
slave_timing[0][32+26].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+26].info_i__max_slave__  = 0.023000000;
slave_timing[0][32+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][32+26].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+26].t_rxd1[0][1] = 1150ns;
slave_timing[0][32+26].t_rxd1[1][0] = 1094ns;
slave_timing[0][32+26].t_rxd1[0][2] = 851ns;
slave_timing[0][32+26].t_rxd1[2][0] = 1383ns;
slave_timing[0][32+26].t_rxd2[0][2] = 1637ns;
slave_timing[0][32+26].t_rxd2[2][0] = 918ns;
slave_timing[0][32+26].t_rxd2[1][2] = 1415ns;
slave_timing[0][32+26].t_rxd2[2][1] = 1186ns;

slave_timing[0][32+27].info_corner          = 2;
slave_timing[0][32+27].info_temp__j__       = 125;
slave_timing[0][32+27].info_i__quite_rec__  = 0.040000000;
slave_timing[0][32+27].info_dtr__ib__       = 1;
slave_timing[0][32+27].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+27].info_i__max_slave__  = 0.025000000;
slave_timing[0][32+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][32+27].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+27].t_rxd1[0][1] = 1100ns;
slave_timing[0][32+27].t_rxd1[1][0] = 1132ns;
slave_timing[0][32+27].t_rxd1[0][2] = 828ns;
slave_timing[0][32+27].t_rxd1[2][0] = 1421ns;
slave_timing[0][32+27].t_rxd2[0][2] = 1503ns;
slave_timing[0][32+27].t_rxd2[2][0] = 981ns;
slave_timing[0][32+27].t_rxd2[1][2] = 1258ns;
slave_timing[0][32+27].t_rxd2[2][1] = 1328ns;

slave_timing[0][32+28].info_corner          = 2;
slave_timing[0][32+28].info_temp__j__       = 125;
slave_timing[0][32+28].info_i__quite_rec__  = 0.040000000;
slave_timing[0][32+28].info_dtr__ib__       = -1;
slave_timing[0][32+28].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+28].info_i__max_slave__  = 0.023000000;
slave_timing[0][32+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][32+28].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+28].t_rxd1[0][1] = 1185ns;
slave_timing[0][32+28].t_rxd1[1][0] = 1186ns;
slave_timing[0][32+28].t_rxd1[0][2] = 921ns;
slave_timing[0][32+28].t_rxd1[2][0] = 1869ns;
slave_timing[0][32+28].t_rxd2[0][2] = 2008ns;
slave_timing[0][32+28].t_rxd2[2][0] = 1413ns;
slave_timing[0][32+28].t_rxd2[1][2] = 1817ns;
slave_timing[0][32+28].t_rxd2[2][1] = 2095ns;

slave_timing[0][32+29].info_corner          = 2;
slave_timing[0][32+29].info_temp__j__       = 125;
slave_timing[0][32+29].info_i__quite_rec__  = 0.040000000;
slave_timing[0][32+29].info_dtr__ib__       = -1;
slave_timing[0][32+29].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+29].info_i__max_slave__  = 0.025000000;
slave_timing[0][32+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][32+29].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+29].t_rxd1[0][1] = 1142ns;
slave_timing[0][32+29].t_rxd1[1][0] = 1212ns;
slave_timing[0][32+29].t_rxd1[0][2] = 901ns;
slave_timing[0][32+29].t_rxd1[2][0] = 1971ns;
slave_timing[0][32+29].t_rxd2[0][2] = 1850ns;
slave_timing[0][32+29].t_rxd2[2][0] = 1534ns;
slave_timing[0][32+29].t_rxd2[1][2] = 1621ns;
slave_timing[0][32+29].t_rxd2[2][1] = 2474ns;

slave_timing[0][32+30].info_corner          = 2;
slave_timing[0][32+30].info_temp__j__       = 125;
slave_timing[0][32+30].info_i__quite_rec__  = 0.040000000;
slave_timing[0][32+30].info_dtr__ib__       = 1;
slave_timing[0][32+30].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+30].info_i__max_slave__  = 0.023000000;
slave_timing[0][32+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][32+30].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+30].t_rxd1[0][1] = 1225ns;
slave_timing[0][32+30].t_rxd1[1][0] = 1146ns;
slave_timing[0][32+30].t_rxd1[0][2] = 939ns;
slave_timing[0][32+30].t_rxd1[2][0] = 1767ns;
slave_timing[0][32+30].t_rxd2[0][2] = 2199ns;
slave_timing[0][32+30].t_rxd2[2][0] = 1297ns;
slave_timing[0][32+30].t_rxd2[1][2] = 2025ns;
slave_timing[0][32+30].t_rxd2[2][1] = 1810ns;

slave_timing[0][32+31].info_corner          = 2;
slave_timing[0][32+31].info_temp__j__       = 125;
slave_timing[0][32+31].info_i__quite_rec__  = 0.040000000;
slave_timing[0][32+31].info_dtr__ib__       = 1;
slave_timing[0][32+31].info_i__offset_rec__ = 0.000000000;
slave_timing[0][32+31].info_i__max_slave__  = 0.025000000;
slave_timing[0][32+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][32+31].info_r__dsi_bus__    = 5.000;

slave_timing[0][32+31].t_rxd1[0][1] = 1178ns;
slave_timing[0][32+31].t_rxd1[1][0] = 1176ns;
slave_timing[0][32+31].t_rxd1[0][2] = 916ns;
slave_timing[0][32+31].t_rxd1[2][0] = 1869ns;
slave_timing[0][32+31].t_rxd2[0][2] = 1979ns;
slave_timing[0][32+31].t_rxd2[2][0] = 1423ns;
slave_timing[0][32+31].t_rxd2[1][2] = 1776ns;
slave_timing[0][32+31].t_rxd2[2][1] = 2136ns;

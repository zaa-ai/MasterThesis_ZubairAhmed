/* ###   interface instances   ###################################################### */

buffer_interrupt_registers_BUF_IRQ_STAT_if buffer_interrupt_registers_BUF_IRQ_STAT (); 
buffer_interrupt_registers_BUF_IRQ_MASK_if buffer_interrupt_registers_BUF_IRQ_MASK (); 
buffer_interrupt_registers_BUF_FILL_WARN_if buffer_interrupt_registers_BUF_FILL_WARN (); 


/* ###   interface instances   ###################################################### */

common_DSI3_block_registers_DSI_ENABLE_if common_DSI3_block_registers_DSI_ENABLE (); 
common_DSI3_block_registers_DSI_CFG_if common_DSI3_block_registers_DSI_CFG (); 
common_DSI3_block_registers_DSI_TX_SHIFT_if common_DSI3_block_registers_DSI_TX_SHIFT (); 
common_DSI3_block_registers_SYNC_IDLE_REG_if common_DSI3_block_registers_SYNC_IDLE_REG (); 
common_DSI3_block_registers_CRM_TIME_if common_DSI3_block_registers_CRM_TIME (); 
common_DSI3_block_registers_CRM_TIME_NR_if common_DSI3_block_registers_CRM_TIME_NR (); 


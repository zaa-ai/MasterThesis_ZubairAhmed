
slave_timing[2][128+0].info_corner          = 1;
slave_timing[2][128+0].info_temp__j__       = -40;
slave_timing[2][128+0].info_i__quite_rec__  = 0.006000000;
slave_timing[2][128+0].info_dtr__ib__       = -1;
slave_timing[2][128+0].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+0].info_i__max_slave__  = 0.023000000;
slave_timing[2][128+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][128+0].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+0].t_rxd1[0][1] = 2144ns;
slave_timing[2][128+0].t_rxd1[1][0] = 2190ns;
slave_timing[2][128+0].t_rxd1[0][2] = 1604ns;
slave_timing[2][128+0].t_rxd1[2][0] = 2653ns;
slave_timing[2][128+0].t_rxd2[0][2] = 2570ns;
slave_timing[2][128+0].t_rxd2[2][0] = 1648ns;
slave_timing[2][128+0].t_rxd2[1][2] = 2118ns;
slave_timing[2][128+0].t_rxd2[2][1] = 2178ns;

slave_timing[2][128+1].info_corner          = 1;
slave_timing[2][128+1].info_temp__j__       = -40;
slave_timing[2][128+1].info_i__quite_rec__  = 0.006000000;
slave_timing[2][128+1].info_dtr__ib__       = -1;
slave_timing[2][128+1].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+1].info_i__max_slave__  = 0.025000000;
slave_timing[2][128+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][128+1].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+1].t_rxd1[0][1] = 2061ns;
slave_timing[2][128+1].t_rxd1[1][0] = 2252ns;
slave_timing[2][128+1].t_rxd1[0][2] = 1573ns;
slave_timing[2][128+1].t_rxd1[2][0] = 2696ns;
slave_timing[2][128+1].t_rxd2[0][2] = 2444ns;
slave_timing[2][128+1].t_rxd2[2][0] = 1756ns;
slave_timing[2][128+1].t_rxd2[1][2] = 1889ns;
slave_timing[2][128+1].t_rxd2[2][1] = 2400ns;

slave_timing[2][128+2].info_corner          = 1;
slave_timing[2][128+2].info_temp__j__       = -40;
slave_timing[2][128+2].info_i__quite_rec__  = 0.006000000;
slave_timing[2][128+2].info_dtr__ib__       = 1;
slave_timing[2][128+2].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+2].info_i__max_slave__  = 0.023000000;
slave_timing[2][128+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][128+2].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+2].t_rxd1[0][1] = 2231ns;
slave_timing[2][128+2].t_rxd1[1][0] = 2117ns;
slave_timing[2][128+2].t_rxd1[0][2] = 1667ns;
slave_timing[2][128+2].t_rxd1[2][0] = 2610ns;
slave_timing[2][128+2].t_rxd2[0][2] = 2749ns;
slave_timing[2][128+2].t_rxd2[2][0] = 1521ns;
slave_timing[2][128+2].t_rxd2[1][2] = 2349ns;
slave_timing[2][128+2].t_rxd2[2][1] = 1977ns;

slave_timing[2][128+3].info_corner          = 1;
slave_timing[2][128+3].info_temp__j__       = -40;
slave_timing[2][128+3].info_i__quite_rec__  = 0.006000000;
slave_timing[2][128+3].info_dtr__ib__       = 1;
slave_timing[2][128+3].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+3].info_i__max_slave__  = 0.025000000;
slave_timing[2][128+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][128+3].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+3].t_rxd1[0][1] = 2136ns;
slave_timing[2][128+3].t_rxd1[1][0] = 2188ns;
slave_timing[2][128+3].t_rxd1[0][2] = 1615ns;
slave_timing[2][128+3].t_rxd1[2][0] = 2653ns;
slave_timing[2][128+3].t_rxd2[0][2] = 2574ns;
slave_timing[2][128+3].t_rxd2[2][0] = 1658ns;
slave_timing[2][128+3].t_rxd2[1][2] = 2103ns;
slave_timing[2][128+3].t_rxd2[2][1] = 2166ns;

slave_timing[2][128+4].info_corner          = 1;
slave_timing[2][128+4].info_temp__j__       = -40;
slave_timing[2][128+4].info_i__quite_rec__  = 0.006000000;
slave_timing[2][128+4].info_dtr__ib__       = -1;
slave_timing[2][128+4].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+4].info_i__max_slave__  = 0.023000000;
slave_timing[2][128+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][128+4].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+4].t_rxd1[0][1] = 2216ns;
slave_timing[2][128+4].t_rxd1[1][0] = 2259ns;
slave_timing[2][128+4].t_rxd1[0][2] = 1668ns;
slave_timing[2][128+4].t_rxd1[2][0] = 2718ns;
slave_timing[2][128+4].t_rxd2[0][2] = 2589ns;
slave_timing[2][128+4].t_rxd2[2][0] = 1661ns;
slave_timing[2][128+4].t_rxd2[1][2] = 2130ns;
slave_timing[2][128+4].t_rxd2[2][1] = 2186ns;

slave_timing[2][128+5].info_corner          = 1;
slave_timing[2][128+5].info_temp__j__       = -40;
slave_timing[2][128+5].info_i__quite_rec__  = 0.006000000;
slave_timing[2][128+5].info_dtr__ib__       = -1;
slave_timing[2][128+5].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+5].info_i__max_slave__  = 0.025000000;
slave_timing[2][128+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][128+5].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+5].t_rxd1[0][1] = 2126ns;
slave_timing[2][128+5].t_rxd1[1][0] = 2320ns;
slave_timing[2][128+5].t_rxd1[0][2] = 1641ns;
slave_timing[2][128+5].t_rxd1[2][0] = 2763ns;
slave_timing[2][128+5].t_rxd2[0][2] = 2464ns;
slave_timing[2][128+5].t_rxd2[2][0] = 1772ns;
slave_timing[2][128+5].t_rxd2[1][2] = 1907ns;
slave_timing[2][128+5].t_rxd2[2][1] = 2420ns;

slave_timing[2][128+6].info_corner          = 1;
slave_timing[2][128+6].info_temp__j__       = -40;
slave_timing[2][128+6].info_i__quite_rec__  = 0.006000000;
slave_timing[2][128+6].info_dtr__ib__       = 1;
slave_timing[2][128+6].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+6].info_i__max_slave__  = 0.023000000;
slave_timing[2][128+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][128+6].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+6].t_rxd1[0][1] = 2295ns;
slave_timing[2][128+6].t_rxd1[1][0] = 2185ns;
slave_timing[2][128+6].t_rxd1[0][2] = 1734ns;
slave_timing[2][128+6].t_rxd1[2][0] = 2678ns;
slave_timing[2][128+6].t_rxd2[0][2] = 2762ns;
slave_timing[2][128+6].t_rxd2[2][0] = 1542ns;
slave_timing[2][128+6].t_rxd2[1][2] = 2360ns;
slave_timing[2][128+6].t_rxd2[2][1] = 1984ns;

slave_timing[2][128+7].info_corner          = 1;
slave_timing[2][128+7].info_temp__j__       = -40;
slave_timing[2][128+7].info_i__quite_rec__  = 0.006000000;
slave_timing[2][128+7].info_dtr__ib__       = 1;
slave_timing[2][128+7].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+7].info_i__max_slave__  = 0.025000000;
slave_timing[2][128+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][128+7].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+7].t_rxd1[0][1] = 2210ns;
slave_timing[2][128+7].t_rxd1[1][0] = 2259ns;
slave_timing[2][128+7].t_rxd1[0][2] = 1680ns;
slave_timing[2][128+7].t_rxd1[2][0] = 2722ns;
slave_timing[2][128+7].t_rxd2[0][2] = 2585ns;
slave_timing[2][128+7].t_rxd2[2][0] = 1676ns;
slave_timing[2][128+7].t_rxd2[1][2] = 2099ns;
slave_timing[2][128+7].t_rxd2[2][1] = 2210ns;

slave_timing[2][128+8].info_corner          = 1;
slave_timing[2][128+8].info_temp__j__       = -40;
slave_timing[2][128+8].info_i__quite_rec__  = 0.003000000;
slave_timing[2][128+8].info_dtr__ib__       = -1;
slave_timing[2][128+8].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+8].info_i__max_slave__  = 0.023000000;
slave_timing[2][128+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][128+8].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+8].t_rxd1[0][1] = 2166ns;
slave_timing[2][128+8].t_rxd1[1][0] = 2170ns;
slave_timing[2][128+8].t_rxd1[0][2] = 1633ns;
slave_timing[2][128+8].t_rxd1[2][0] = 2636ns;
slave_timing[2][128+8].t_rxd2[0][2] = 2607ns;
slave_timing[2][128+8].t_rxd2[2][0] = 1638ns;
slave_timing[2][128+8].t_rxd2[1][2] = 2143ns;
slave_timing[2][128+8].t_rxd2[2][1] = 2161ns;

slave_timing[2][128+9].info_corner          = 1;
slave_timing[2][128+9].info_temp__j__       = -40;
slave_timing[2][128+9].info_i__quite_rec__  = 0.003000000;
slave_timing[2][128+9].info_dtr__ib__       = -1;
slave_timing[2][128+9].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+9].info_i__max_slave__  = 0.025000000;
slave_timing[2][128+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][128+9].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+9].t_rxd1[0][1] = 2081ns;
slave_timing[2][128+9].t_rxd1[1][0] = 2226ns;
slave_timing[2][128+9].t_rxd1[0][2] = 1586ns;
slave_timing[2][128+9].t_rxd1[2][0] = 2682ns;
slave_timing[2][128+9].t_rxd2[0][2] = 2457ns;
slave_timing[2][128+9].t_rxd2[2][0] = 1751ns;
slave_timing[2][128+9].t_rxd2[1][2] = 1907ns;
slave_timing[2][128+9].t_rxd2[2][1] = 2390ns;

slave_timing[2][128+10].info_corner          = 1;
slave_timing[2][128+10].info_temp__j__       = -40;
slave_timing[2][128+10].info_i__quite_rec__  = 0.003000000;
slave_timing[2][128+10].info_dtr__ib__       = 1;
slave_timing[2][128+10].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+10].info_i__max_slave__  = 0.023000000;
slave_timing[2][128+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][128+10].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+10].t_rxd1[0][1] = 2243ns;
slave_timing[2][128+10].t_rxd1[1][0] = 2093ns;
slave_timing[2][128+10].t_rxd1[0][2] = 1677ns;
slave_timing[2][128+10].t_rxd1[2][0] = 2592ns;
slave_timing[2][128+10].t_rxd2[0][2] = 2767ns;
slave_timing[2][128+10].t_rxd2[2][0] = 1517ns;
slave_timing[2][128+10].t_rxd2[1][2] = 2372ns;
slave_timing[2][128+10].t_rxd2[2][1] = 1956ns;

slave_timing[2][128+11].info_corner          = 1;
slave_timing[2][128+11].info_temp__j__       = -40;
slave_timing[2][128+11].info_i__quite_rec__  = 0.003000000;
slave_timing[2][128+11].info_dtr__ib__       = 1;
slave_timing[2][128+11].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+11].info_i__max_slave__  = 0.025000000;
slave_timing[2][128+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][128+11].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+11].t_rxd1[0][1] = 2158ns;
slave_timing[2][128+11].t_rxd1[1][0] = 2159ns;
slave_timing[2][128+11].t_rxd1[0][2] = 1627ns;
slave_timing[2][128+11].t_rxd1[2][0] = 2640ns;
slave_timing[2][128+11].t_rxd2[0][2] = 2588ns;
slave_timing[2][128+11].t_rxd2[2][0] = 1650ns;
slave_timing[2][128+11].t_rxd2[1][2] = 2105ns;
slave_timing[2][128+11].t_rxd2[2][1] = 2190ns;

slave_timing[2][128+12].info_corner          = 1;
slave_timing[2][128+12].info_temp__j__       = -40;
slave_timing[2][128+12].info_i__quite_rec__  = 0.003000000;
slave_timing[2][128+12].info_dtr__ib__       = -1;
slave_timing[2][128+12].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+12].info_i__max_slave__  = 0.023000000;
slave_timing[2][128+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][128+12].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+12].t_rxd1[0][1] = 2240ns;
slave_timing[2][128+12].t_rxd1[1][0] = 2237ns;
slave_timing[2][128+12].t_rxd1[0][2] = 1701ns;
slave_timing[2][128+12].t_rxd1[2][0] = 2709ns;
slave_timing[2][128+12].t_rxd2[0][2] = 2622ns;
slave_timing[2][128+12].t_rxd2[2][0] = 1651ns;
slave_timing[2][128+12].t_rxd2[1][2] = 2153ns;
slave_timing[2][128+12].t_rxd2[2][1] = 2176ns;

slave_timing[2][128+13].info_corner          = 1;
slave_timing[2][128+13].info_temp__j__       = -40;
slave_timing[2][128+13].info_i__quite_rec__  = 0.003000000;
slave_timing[2][128+13].info_dtr__ib__       = -1;
slave_timing[2][128+13].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+13].info_i__max_slave__  = 0.025000000;
slave_timing[2][128+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][128+13].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+13].t_rxd1[0][1] = 2157ns;
slave_timing[2][128+13].t_rxd1[1][0] = 2306ns;
slave_timing[2][128+13].t_rxd1[0][2] = 1654ns;
slave_timing[2][128+13].t_rxd1[2][0] = 2750ns;
slave_timing[2][128+13].t_rxd2[0][2] = 2475ns;
slave_timing[2][128+13].t_rxd2[2][0] = 1766ns;
slave_timing[2][128+13].t_rxd2[1][2] = 1930ns;
slave_timing[2][128+13].t_rxd2[2][1] = 2408ns;

slave_timing[2][128+14].info_corner          = 1;
slave_timing[2][128+14].info_temp__j__       = -40;
slave_timing[2][128+14].info_i__quite_rec__  = 0.003000000;
slave_timing[2][128+14].info_dtr__ib__       = 1;
slave_timing[2][128+14].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+14].info_i__max_slave__  = 0.023000000;
slave_timing[2][128+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][128+14].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+14].t_rxd1[0][1] = 2323ns;
slave_timing[2][128+14].t_rxd1[1][0] = 2163ns;
slave_timing[2][128+14].t_rxd1[0][2] = 1745ns;
slave_timing[2][128+14].t_rxd1[2][0] = 2660ns;
slave_timing[2][128+14].t_rxd2[0][2] = 2777ns;
slave_timing[2][128+14].t_rxd2[2][0] = 1536ns;
slave_timing[2][128+14].t_rxd2[1][2] = 2380ns;
slave_timing[2][128+14].t_rxd2[2][1] = 1962ns;

slave_timing[2][128+15].info_corner          = 1;
slave_timing[2][128+15].info_temp__j__       = -40;
slave_timing[2][128+15].info_i__quite_rec__  = 0.003000000;
slave_timing[2][128+15].info_dtr__ib__       = 1;
slave_timing[2][128+15].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+15].info_i__max_slave__  = 0.025000000;
slave_timing[2][128+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][128+15].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+15].t_rxd1[0][1] = 2232ns;
slave_timing[2][128+15].t_rxd1[1][0] = 2230ns;
slave_timing[2][128+15].t_rxd1[0][2] = 1694ns;
slave_timing[2][128+15].t_rxd1[2][0] = 2706ns;
slave_timing[2][128+15].t_rxd2[0][2] = 2600ns;
slave_timing[2][128+15].t_rxd2[2][0] = 1664ns;
slave_timing[2][128+15].t_rxd2[1][2] = 2118ns;
slave_timing[2][128+15].t_rxd2[2][1] = 2200ns;

slave_timing[2][128+16].info_corner          = 1;
slave_timing[2][128+16].info_temp__j__       = -40;
slave_timing[2][128+16].info_i__quite_rec__  = 0.000000000;
slave_timing[2][128+16].info_dtr__ib__       = -1;
slave_timing[2][128+16].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+16].info_i__max_slave__  = 0.023000000;
slave_timing[2][128+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][128+16].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+16].t_rxd1[0][1] = 2146ns;
slave_timing[2][128+16].t_rxd1[1][0] = 2168ns;
slave_timing[2][128+16].t_rxd1[0][2] = 1623ns;
slave_timing[2][128+16].t_rxd1[2][0] = 2647ns;
slave_timing[2][128+16].t_rxd2[0][2] = 2597ns;
slave_timing[2][128+16].t_rxd2[2][0] = 1644ns;
slave_timing[2][128+16].t_rxd2[1][2] = 2122ns;
slave_timing[2][128+16].t_rxd2[2][1] = 2181ns;

slave_timing[2][128+17].info_corner          = 1;
slave_timing[2][128+17].info_temp__j__       = -40;
slave_timing[2][128+17].info_i__quite_rec__  = 0.000000000;
slave_timing[2][128+17].info_dtr__ib__       = -1;
slave_timing[2][128+17].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+17].info_i__max_slave__  = 0.025000000;
slave_timing[2][128+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][128+17].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+17].t_rxd1[0][1] = 2063ns;
slave_timing[2][128+17].t_rxd1[1][0] = 2237ns;
slave_timing[2][128+17].t_rxd1[0][2] = 1578ns;
slave_timing[2][128+17].t_rxd1[2][0] = 2692ns;
slave_timing[2][128+17].t_rxd2[0][2] = 2453ns;
slave_timing[2][128+17].t_rxd2[2][0] = 1759ns;
slave_timing[2][128+17].t_rxd2[1][2] = 1899ns;
slave_timing[2][128+17].t_rxd2[2][1] = 2407ns;

slave_timing[2][128+18].info_corner          = 1;
slave_timing[2][128+18].info_temp__j__       = -40;
slave_timing[2][128+18].info_i__quite_rec__  = 0.000000000;
slave_timing[2][128+18].info_dtr__ib__       = 1;
slave_timing[2][128+18].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+18].info_i__max_slave__  = 0.023000000;
slave_timing[2][128+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][128+18].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+18].t_rxd1[0][1] = 2219ns;
slave_timing[2][128+18].t_rxd1[1][0] = 2105ns;
slave_timing[2][128+18].t_rxd1[0][2] = 1665ns;
slave_timing[2][128+18].t_rxd1[2][0] = 2604ns;
slave_timing[2][128+18].t_rxd2[0][2] = 2752ns;
slave_timing[2][128+18].t_rxd2[2][0] = 1516ns;
slave_timing[2][128+18].t_rxd2[1][2] = 2352ns;
slave_timing[2][128+18].t_rxd2[2][1] = 1960ns;

slave_timing[2][128+19].info_corner          = 1;
slave_timing[2][128+19].info_temp__j__       = -40;
slave_timing[2][128+19].info_i__quite_rec__  = 0.000000000;
slave_timing[2][128+19].info_dtr__ib__       = 1;
slave_timing[2][128+19].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+19].info_i__max_slave__  = 0.025000000;
slave_timing[2][128+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][128+19].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+19].t_rxd1[0][1] = 2142ns;
slave_timing[2][128+19].t_rxd1[1][0] = 2180ns;
slave_timing[2][128+19].t_rxd1[0][2] = 1618ns;
slave_timing[2][128+19].t_rxd1[2][0] = 2651ns;
slave_timing[2][128+19].t_rxd2[0][2] = 2568ns;
slave_timing[2][128+19].t_rxd2[2][0] = 1655ns;
slave_timing[2][128+19].t_rxd2[1][2] = 2081ns;
slave_timing[2][128+19].t_rxd2[2][1] = 2196ns;

slave_timing[2][128+20].info_corner          = 1;
slave_timing[2][128+20].info_temp__j__       = -40;
slave_timing[2][128+20].info_i__quite_rec__  = 0.000000000;
slave_timing[2][128+20].info_dtr__ib__       = -1;
slave_timing[2][128+20].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+20].info_i__max_slave__  = 0.023000000;
slave_timing[2][128+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][128+20].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+20].t_rxd1[0][1] = 2214ns;
slave_timing[2][128+20].t_rxd1[1][0] = 2238ns;
slave_timing[2][128+20].t_rxd1[0][2] = 1693ns;
slave_timing[2][128+20].t_rxd1[2][0] = 2715ns;
slave_timing[2][128+20].t_rxd2[0][2] = 2608ns;
slave_timing[2][128+20].t_rxd2[2][0] = 1662ns;
slave_timing[2][128+20].t_rxd2[1][2] = 2127ns;
slave_timing[2][128+20].t_rxd2[2][1] = 2193ns;

slave_timing[2][128+21].info_corner          = 1;
slave_timing[2][128+21].info_temp__j__       = -40;
slave_timing[2][128+21].info_i__quite_rec__  = 0.000000000;
slave_timing[2][128+21].info_dtr__ib__       = -1;
slave_timing[2][128+21].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+21].info_i__max_slave__  = 0.025000000;
slave_timing[2][128+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][128+21].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+21].t_rxd1[0][1] = 2144ns;
slave_timing[2][128+21].t_rxd1[1][0] = 2305ns;
slave_timing[2][128+21].t_rxd1[0][2] = 1645ns;
slave_timing[2][128+21].t_rxd1[2][0] = 2757ns;
slave_timing[2][128+21].t_rxd2[0][2] = 2466ns;
slave_timing[2][128+21].t_rxd2[2][0] = 1774ns;
slave_timing[2][128+21].t_rxd2[1][2] = 1944ns;
slave_timing[2][128+21].t_rxd2[2][1] = 2382ns;

slave_timing[2][128+22].info_corner          = 1;
slave_timing[2][128+22].info_temp__j__       = -40;
slave_timing[2][128+22].info_i__quite_rec__  = 0.000000000;
slave_timing[2][128+22].info_dtr__ib__       = 1;
slave_timing[2][128+22].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+22].info_i__max_slave__  = 0.023000000;
slave_timing[2][128+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][128+22].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+22].t_rxd1[0][1] = 2291ns;
slave_timing[2][128+22].t_rxd1[1][0] = 2189ns;
slave_timing[2][128+22].t_rxd1[0][2] = 1735ns;
slave_timing[2][128+22].t_rxd1[2][0] = 2673ns;
slave_timing[2][128+22].t_rxd2[0][2] = 2758ns;
slave_timing[2][128+22].t_rxd2[2][0] = 1539ns;
slave_timing[2][128+22].t_rxd2[1][2] = 2365ns;
slave_timing[2][128+22].t_rxd2[2][1] = 1974ns;

slave_timing[2][128+23].info_corner          = 1;
slave_timing[2][128+23].info_temp__j__       = -40;
slave_timing[2][128+23].info_i__quite_rec__  = 0.000000000;
slave_timing[2][128+23].info_dtr__ib__       = 1;
slave_timing[2][128+23].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+23].info_i__max_slave__  = 0.025000000;
slave_timing[2][128+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][128+23].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+23].t_rxd1[0][1] = 2212ns;
slave_timing[2][128+23].t_rxd1[1][0] = 2251ns;
slave_timing[2][128+23].t_rxd1[0][2] = 1682ns;
slave_timing[2][128+23].t_rxd1[2][0] = 2717ns;
slave_timing[2][128+23].t_rxd2[0][2] = 2586ns;
slave_timing[2][128+23].t_rxd2[2][0] = 1666ns;
slave_timing[2][128+23].t_rxd2[1][2] = 2100ns;
slave_timing[2][128+23].t_rxd2[2][1] = 2177ns;

slave_timing[2][128+24].info_corner          = 1;
slave_timing[2][128+24].info_temp__j__       = -40;
slave_timing[2][128+24].info_i__quite_rec__  = 0.040000000;
slave_timing[2][128+24].info_dtr__ib__       = -1;
slave_timing[2][128+24].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+24].info_i__max_slave__  = 0.023000000;
slave_timing[2][128+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][128+24].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+24].t_rxd1[0][1] = 2167ns;
slave_timing[2][128+24].t_rxd1[1][0] = 2146ns;
slave_timing[2][128+24].t_rxd1[0][2] = 1628ns;
slave_timing[2][128+24].t_rxd1[2][0] = 2625ns;
slave_timing[2][128+24].t_rxd2[0][2] = 2612ns;
slave_timing[2][128+24].t_rxd2[2][0] = 1635ns;
slave_timing[2][128+24].t_rxd2[1][2] = 2136ns;
slave_timing[2][128+24].t_rxd2[2][1] = 2155ns;

slave_timing[2][128+25].info_corner          = 1;
slave_timing[2][128+25].info_temp__j__       = -40;
slave_timing[2][128+25].info_i__quite_rec__  = 0.040000000;
slave_timing[2][128+25].info_dtr__ib__       = -1;
slave_timing[2][128+25].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+25].info_i__max_slave__  = 0.025000000;
slave_timing[2][128+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][128+25].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+25].t_rxd1[0][1] = 2080ns;
slave_timing[2][128+25].t_rxd1[1][0] = 2218ns;
slave_timing[2][128+25].t_rxd1[0][2] = 1581ns;
slave_timing[2][128+25].t_rxd1[2][0] = 2670ns;
slave_timing[2][128+25].t_rxd2[0][2] = 2466ns;
slave_timing[2][128+25].t_rxd2[2][0] = 1748ns;
slave_timing[2][128+25].t_rxd2[1][2] = 1907ns;
slave_timing[2][128+25].t_rxd2[2][1] = 2390ns;

slave_timing[2][128+26].info_corner          = 1;
slave_timing[2][128+26].info_temp__j__       = -40;
slave_timing[2][128+26].info_i__quite_rec__  = 0.040000000;
slave_timing[2][128+26].info_dtr__ib__       = 1;
slave_timing[2][128+26].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+26].info_i__max_slave__  = 0.023000000;
slave_timing[2][128+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][128+26].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+26].t_rxd1[0][1] = 2213ns;
slave_timing[2][128+26].t_rxd1[1][0] = 2118ns;
slave_timing[2][128+26].t_rxd1[0][2] = 1659ns;
slave_timing[2][128+26].t_rxd1[2][0] = 2600ns;
slave_timing[2][128+26].t_rxd2[0][2] = 2748ns;
slave_timing[2][128+26].t_rxd2[2][0] = 1533ns;
slave_timing[2][128+26].t_rxd2[1][2] = 2344ns;
slave_timing[2][128+26].t_rxd2[2][1] = 1973ns;

slave_timing[2][128+27].info_corner          = 1;
slave_timing[2][128+27].info_temp__j__       = -40;
slave_timing[2][128+27].info_i__quite_rec__  = 0.040000000;
slave_timing[2][128+27].info_dtr__ib__       = 1;
slave_timing[2][128+27].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+27].info_i__max_slave__  = 0.025000000;
slave_timing[2][128+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][128+27].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+27].t_rxd1[0][1] = 2135ns;
slave_timing[2][128+27].t_rxd1[1][0] = 2188ns;
slave_timing[2][128+27].t_rxd1[0][2] = 1609ns;
slave_timing[2][128+27].t_rxd1[2][0] = 2645ns;
slave_timing[2][128+27].t_rxd2[0][2] = 2566ns;
slave_timing[2][128+27].t_rxd2[2][0] = 1664ns;
slave_timing[2][128+27].t_rxd2[1][2] = 2087ns;
slave_timing[2][128+27].t_rxd2[2][1] = 2182ns;

slave_timing[2][128+28].info_corner          = 1;
slave_timing[2][128+28].info_temp__j__       = -40;
slave_timing[2][128+28].info_i__quite_rec__  = 0.040000000;
slave_timing[2][128+28].info_dtr__ib__       = -1;
slave_timing[2][128+28].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+28].info_i__max_slave__  = 0.023000000;
slave_timing[2][128+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][128+28].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+28].t_rxd1[0][1] = 2193ns;
slave_timing[2][128+28].t_rxd1[1][0] = 2194ns;
slave_timing[2][128+28].t_rxd1[0][2] = 1668ns;
slave_timing[2][128+28].t_rxd1[2][0] = 2668ns;
slave_timing[2][128+28].t_rxd2[0][2] = 2616ns;
slave_timing[2][128+28].t_rxd2[2][0] = 1648ns;
slave_timing[2][128+28].t_rxd2[1][2] = 2147ns;
slave_timing[2][128+28].t_rxd2[2][1] = 2133ns;

slave_timing[2][128+29].info_corner          = 1;
slave_timing[2][128+29].info_temp__j__       = -40;
slave_timing[2][128+29].info_i__quite_rec__  = 0.040000000;
slave_timing[2][128+29].info_dtr__ib__       = -1;
slave_timing[2][128+29].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+29].info_i__max_slave__  = 0.025000000;
slave_timing[2][128+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][128+29].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+29].t_rxd1[0][1] = 2113ns;
slave_timing[2][128+29].t_rxd1[1][0] = 2261ns;
slave_timing[2][128+29].t_rxd1[0][2] = 1602ns;
slave_timing[2][128+29].t_rxd1[2][0] = 2715ns;
slave_timing[2][128+29].t_rxd2[0][2] = 2455ns;
slave_timing[2][128+29].t_rxd2[2][0] = 1764ns;
slave_timing[2][128+29].t_rxd2[1][2] = 1920ns;
slave_timing[2][128+29].t_rxd2[2][1] = 2396ns;

slave_timing[2][128+30].info_corner          = 1;
slave_timing[2][128+30].info_temp__j__       = -40;
slave_timing[2][128+30].info_i__quite_rec__  = 0.040000000;
slave_timing[2][128+30].info_dtr__ib__       = 1;
slave_timing[2][128+30].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+30].info_i__max_slave__  = 0.023000000;
slave_timing[2][128+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][128+30].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+30].t_rxd1[0][1] = 2259ns;
slave_timing[2][128+30].t_rxd1[1][0] = 2163ns;
slave_timing[2][128+30].t_rxd1[0][2] = 1698ns;
slave_timing[2][128+30].t_rxd1[2][0] = 2645ns;
slave_timing[2][128+30].t_rxd2[0][2] = 2756ns;
slave_timing[2][128+30].t_rxd2[2][0] = 1548ns;
slave_timing[2][128+30].t_rxd2[1][2] = 2350ns;
slave_timing[2][128+30].t_rxd2[2][1] = 1993ns;

slave_timing[2][128+31].info_corner          = 1;
slave_timing[2][128+31].info_temp__j__       = -40;
slave_timing[2][128+31].info_i__quite_rec__  = 0.040000000;
slave_timing[2][128+31].info_dtr__ib__       = 1;
slave_timing[2][128+31].info_i__offset_rec__ = 0.000000000;
slave_timing[2][128+31].info_i__max_slave__  = 0.025000000;
slave_timing[2][128+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][128+31].info_r__dsi_bus__    = 5.000;

slave_timing[2][128+31].t_rxd1[0][1] = 2162ns;
slave_timing[2][128+31].t_rxd1[1][0] = 2221ns;
slave_timing[2][128+31].t_rxd1[0][2] = 1649ns;
slave_timing[2][128+31].t_rxd1[2][0] = 2686ns;
slave_timing[2][128+31].t_rxd2[0][2] = 2584ns;
slave_timing[2][128+31].t_rxd2[2][0] = 1679ns;
slave_timing[2][128+31].t_rxd2[1][2] = 2103ns;
slave_timing[2][128+31].t_rxd2[2][1] = 2225ns;

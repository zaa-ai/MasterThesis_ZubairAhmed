import dsi3_master_pkg::*;

`include "slave_rxd_timing.svh"
`include "slave_timing_container.svh"
`include "dsi3_chip_distribution.svh"

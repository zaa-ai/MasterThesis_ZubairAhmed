
slave_timing[2][192+0].info_corner          = 3;
slave_timing[2][192+0].info_temp__j__       = -40;
slave_timing[2][192+0].info_i__quite_rec__  = 0.006000000;
slave_timing[2][192+0].info_dtr__ib__       = -1;
slave_timing[2][192+0].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+0].info_i__max_slave__  = 0.023000000;
slave_timing[2][192+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][192+0].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+0].t_rxd1[0][1] = 2176ns;
slave_timing[2][192+0].t_rxd1[1][0] = 2216ns;
slave_timing[2][192+0].t_rxd1[0][2] = 1648ns;
slave_timing[2][192+0].t_rxd1[2][0] = 2687ns;
slave_timing[2][192+0].t_rxd2[0][2] = 2634ns;
slave_timing[2][192+0].t_rxd2[2][0] = 1674ns;
slave_timing[2][192+0].t_rxd2[1][2] = 2146ns;
slave_timing[2][192+0].t_rxd2[2][1] = 2221ns;

slave_timing[2][192+1].info_corner          = 3;
slave_timing[2][192+1].info_temp__j__       = -40;
slave_timing[2][192+1].info_i__quite_rec__  = 0.006000000;
slave_timing[2][192+1].info_dtr__ib__       = -1;
slave_timing[2][192+1].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+1].info_i__max_slave__  = 0.025000000;
slave_timing[2][192+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][192+1].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+1].t_rxd1[0][1] = 2095ns;
slave_timing[2][192+1].t_rxd1[1][0] = 2283ns;
slave_timing[2][192+1].t_rxd1[0][2] = 1601ns;
slave_timing[2][192+1].t_rxd1[2][0] = 2740ns;
slave_timing[2][192+1].t_rxd2[0][2] = 2489ns;
slave_timing[2][192+1].t_rxd2[2][0] = 1788ns;
slave_timing[2][192+1].t_rxd2[1][2] = 1916ns;
slave_timing[2][192+1].t_rxd2[2][1] = 2443ns;

slave_timing[2][192+2].info_corner          = 3;
slave_timing[2][192+2].info_temp__j__       = -40;
slave_timing[2][192+2].info_i__quite_rec__  = 0.006000000;
slave_timing[2][192+2].info_dtr__ib__       = 1;
slave_timing[2][192+2].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+2].info_i__max_slave__  = 0.023000000;
slave_timing[2][192+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][192+2].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+2].t_rxd1[0][1] = 2238ns;
slave_timing[2][192+2].t_rxd1[1][0] = 2161ns;
slave_timing[2][192+2].t_rxd1[0][2] = 1673ns;
slave_timing[2][192+2].t_rxd1[2][0] = 2650ns;
slave_timing[2][192+2].t_rxd2[0][2] = 2764ns;
slave_timing[2][192+2].t_rxd2[2][0] = 1559ns;
slave_timing[2][192+2].t_rxd2[1][2] = 2342ns;
slave_timing[2][192+2].t_rxd2[2][1] = 2040ns;

slave_timing[2][192+3].info_corner          = 3;
slave_timing[2][192+3].info_temp__j__       = -40;
slave_timing[2][192+3].info_i__quite_rec__  = 0.006000000;
slave_timing[2][192+3].info_dtr__ib__       = 1;
slave_timing[2][192+3].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+3].info_i__max_slave__  = 0.025000000;
slave_timing[2][192+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][192+3].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+3].t_rxd1[0][1] = 2153ns;
slave_timing[2][192+3].t_rxd1[1][0] = 2231ns;
slave_timing[2][192+3].t_rxd1[0][2] = 1636ns;
slave_timing[2][192+3].t_rxd1[2][0] = 2704ns;
slave_timing[2][192+3].t_rxd2[0][2] = 2592ns;
slave_timing[2][192+3].t_rxd2[2][0] = 1705ns;
slave_timing[2][192+3].t_rxd2[1][2] = 2122ns;
slave_timing[2][192+3].t_rxd2[2][1] = 2255ns;

slave_timing[2][192+4].info_corner          = 3;
slave_timing[2][192+4].info_temp__j__       = -40;
slave_timing[2][192+4].info_i__quite_rec__  = 0.006000000;
slave_timing[2][192+4].info_dtr__ib__       = -1;
slave_timing[2][192+4].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+4].info_i__max_slave__  = 0.023000000;
slave_timing[2][192+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][192+4].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+4].t_rxd1[0][1] = 2257ns;
slave_timing[2][192+4].t_rxd1[1][0] = 2294ns;
slave_timing[2][192+4].t_rxd1[0][2] = 1723ns;
slave_timing[2][192+4].t_rxd1[2][0] = 2762ns;
slave_timing[2][192+4].t_rxd2[0][2] = 2652ns;
slave_timing[2][192+4].t_rxd2[2][0] = 1688ns;
slave_timing[2][192+4].t_rxd2[1][2] = 2162ns;
slave_timing[2][192+4].t_rxd2[2][1] = 2236ns;

slave_timing[2][192+5].info_corner          = 3;
slave_timing[2][192+5].info_temp__j__       = -40;
slave_timing[2][192+5].info_i__quite_rec__  = 0.006000000;
slave_timing[2][192+5].info_dtr__ib__       = -1;
slave_timing[2][192+5].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+5].info_i__max_slave__  = 0.025000000;
slave_timing[2][192+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][192+5].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+5].t_rxd1[0][1] = 2170ns;
slave_timing[2][192+5].t_rxd1[1][0] = 2355ns;
slave_timing[2][192+5].t_rxd1[0][2] = 1669ns;
slave_timing[2][192+5].t_rxd1[2][0] = 2811ns;
slave_timing[2][192+5].t_rxd2[0][2] = 2508ns;
slave_timing[2][192+5].t_rxd2[2][0] = 1808ns;
slave_timing[2][192+5].t_rxd2[1][2] = 1929ns;
slave_timing[2][192+5].t_rxd2[2][1] = 2464ns;

slave_timing[2][192+6].info_corner          = 3;
slave_timing[2][192+6].info_temp__j__       = -40;
slave_timing[2][192+6].info_i__quite_rec__  = 0.006000000;
slave_timing[2][192+6].info_dtr__ib__       = 1;
slave_timing[2][192+6].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+6].info_i__max_slave__  = 0.023000000;
slave_timing[2][192+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][192+6].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+6].t_rxd1[0][1] = 2314ns;
slave_timing[2][192+6].t_rxd1[1][0] = 2235ns;
slave_timing[2][192+6].t_rxd1[0][2] = 1749ns;
slave_timing[2][192+6].t_rxd1[2][0] = 2723ns;
slave_timing[2][192+6].t_rxd2[0][2] = 2782ns;
slave_timing[2][192+6].t_rxd2[2][0] = 1575ns;
slave_timing[2][192+6].t_rxd2[1][2] = 2344ns;
slave_timing[2][192+6].t_rxd2[2][1] = 2052ns;

slave_timing[2][192+7].info_corner          = 3;
slave_timing[2][192+7].info_temp__j__       = -40;
slave_timing[2][192+7].info_i__quite_rec__  = 0.006000000;
slave_timing[2][192+7].info_dtr__ib__       = 1;
slave_timing[2][192+7].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+7].info_i__max_slave__  = 0.025000000;
slave_timing[2][192+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][192+7].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+7].t_rxd1[0][1] = 2228ns;
slave_timing[2][192+7].t_rxd1[1][0] = 2303ns;
slave_timing[2][192+7].t_rxd1[0][2] = 1700ns;
slave_timing[2][192+7].t_rxd1[2][0] = 2775ns;
slave_timing[2][192+7].t_rxd2[0][2] = 2609ns;
slave_timing[2][192+7].t_rxd2[2][0] = 1719ns;
slave_timing[2][192+7].t_rxd2[1][2] = 2097ns;
slave_timing[2][192+7].t_rxd2[2][1] = 2291ns;

slave_timing[2][192+8].info_corner          = 3;
slave_timing[2][192+8].info_temp__j__       = -40;
slave_timing[2][192+8].info_i__quite_rec__  = 0.003000000;
slave_timing[2][192+8].info_dtr__ib__       = -1;
slave_timing[2][192+8].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+8].info_i__max_slave__  = 0.023000000;
slave_timing[2][192+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][192+8].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+8].t_rxd1[0][1] = 2177ns;
slave_timing[2][192+8].t_rxd1[1][0] = 2234ns;
slave_timing[2][192+8].t_rxd1[0][2] = 1641ns;
slave_timing[2][192+8].t_rxd1[2][0] = 2703ns;
slave_timing[2][192+8].t_rxd2[0][2] = 2627ns;
slave_timing[2][192+8].t_rxd2[2][0] = 1676ns;
slave_timing[2][192+8].t_rxd2[1][2] = 2164ns;
slave_timing[2][192+8].t_rxd2[2][1] = 2191ns;

slave_timing[2][192+9].info_corner          = 3;
slave_timing[2][192+9].info_temp__j__       = -40;
slave_timing[2][192+9].info_i__quite_rec__  = 0.003000000;
slave_timing[2][192+9].info_dtr__ib__       = -1;
slave_timing[2][192+9].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+9].info_i__max_slave__  = 0.025000000;
slave_timing[2][192+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][192+9].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+9].t_rxd1[0][1] = 2089ns;
slave_timing[2][192+9].t_rxd1[1][0] = 2295ns;
slave_timing[2][192+9].t_rxd1[0][2] = 1599ns;
slave_timing[2][192+9].t_rxd1[2][0] = 2752ns;
slave_timing[2][192+9].t_rxd2[0][2] = 2481ns;
slave_timing[2][192+9].t_rxd2[2][0] = 1792ns;
slave_timing[2][192+9].t_rxd2[1][2] = 1907ns;
slave_timing[2][192+9].t_rxd2[2][1] = 2462ns;

slave_timing[2][192+10].info_corner          = 3;
slave_timing[2][192+10].info_temp__j__       = -40;
slave_timing[2][192+10].info_i__quite_rec__  = 0.003000000;
slave_timing[2][192+10].info_dtr__ib__       = 1;
slave_timing[2][192+10].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+10].info_i__max_slave__  = 0.023000000;
slave_timing[2][192+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][192+10].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+10].t_rxd1[0][1] = 2237ns;
slave_timing[2][192+10].t_rxd1[1][0] = 2169ns;
slave_timing[2][192+10].t_rxd1[0][2] = 1674ns;
slave_timing[2][192+10].t_rxd1[2][0] = 2670ns;
slave_timing[2][192+10].t_rxd2[0][2] = 2757ns;
slave_timing[2][192+10].t_rxd2[2][0] = 1580ns;
slave_timing[2][192+10].t_rxd2[1][2] = 2332ns;
slave_timing[2][192+10].t_rxd2[2][1] = 2056ns;

slave_timing[2][192+11].info_corner          = 3;
slave_timing[2][192+11].info_temp__j__       = -40;
slave_timing[2][192+11].info_i__quite_rec__  = 0.003000000;
slave_timing[2][192+11].info_dtr__ib__       = 1;
slave_timing[2][192+11].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+11].info_i__max_slave__  = 0.025000000;
slave_timing[2][192+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][192+11].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+11].t_rxd1[0][1] = 2149ns;
slave_timing[2][192+11].t_rxd1[1][0] = 2227ns;
slave_timing[2][192+11].t_rxd1[0][2] = 1632ns;
slave_timing[2][192+11].t_rxd1[2][0] = 2710ns;
slave_timing[2][192+11].t_rxd2[0][2] = 2589ns;
slave_timing[2][192+11].t_rxd2[2][0] = 1708ns;
slave_timing[2][192+11].t_rxd2[1][2] = 2081ns;
slave_timing[2][192+11].t_rxd2[2][1] = 2277ns;

slave_timing[2][192+12].info_corner          = 3;
slave_timing[2][192+12].info_temp__j__       = -40;
slave_timing[2][192+12].info_i__quite_rec__  = 0.003000000;
slave_timing[2][192+12].info_dtr__ib__       = -1;
slave_timing[2][192+12].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+12].info_i__max_slave__  = 0.023000000;
slave_timing[2][192+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][192+12].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+12].t_rxd1[0][1] = 2289ns;
slave_timing[2][192+12].t_rxd1[1][0] = 2275ns;
slave_timing[2][192+12].t_rxd1[0][2] = 1715ns;
slave_timing[2][192+12].t_rxd1[2][0] = 2780ns;
slave_timing[2][192+12].t_rxd2[0][2] = 2643ns;
slave_timing[2][192+12].t_rxd2[2][0] = 1697ns;
slave_timing[2][192+12].t_rxd2[1][2] = 2178ns;
slave_timing[2][192+12].t_rxd2[2][1] = 2215ns;

slave_timing[2][192+13].info_corner          = 3;
slave_timing[2][192+13].info_temp__j__       = -40;
slave_timing[2][192+13].info_i__quite_rec__  = 0.003000000;
slave_timing[2][192+13].info_dtr__ib__       = -1;
slave_timing[2][192+13].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+13].info_i__max_slave__  = 0.025000000;
slave_timing[2][192+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][192+13].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+13].t_rxd1[0][1] = 2173ns;
slave_timing[2][192+13].t_rxd1[1][0] = 2378ns;
slave_timing[2][192+13].t_rxd1[0][2] = 1673ns;
slave_timing[2][192+13].t_rxd1[2][0] = 2821ns;
slave_timing[2][192+13].t_rxd2[0][2] = 2502ns;
slave_timing[2][192+13].t_rxd2[2][0] = 1808ns;
slave_timing[2][192+13].t_rxd2[1][2] = 1925ns;
slave_timing[2][192+13].t_rxd2[2][1] = 2473ns;

slave_timing[2][192+14].info_corner          = 3;
slave_timing[2][192+14].info_temp__j__       = -40;
slave_timing[2][192+14].info_i__quite_rec__  = 0.003000000;
slave_timing[2][192+14].info_dtr__ib__       = 1;
slave_timing[2][192+14].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+14].info_i__max_slave__  = 0.023000000;
slave_timing[2][192+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][192+14].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+14].t_rxd1[0][1] = 2309ns;
slave_timing[2][192+14].t_rxd1[1][0] = 2243ns;
slave_timing[2][192+14].t_rxd1[0][2] = 1749ns;
slave_timing[2][192+14].t_rxd1[2][0] = 2731ns;
slave_timing[2][192+14].t_rxd2[0][2] = 2779ns;
slave_timing[2][192+14].t_rxd2[2][0] = 1594ns;
slave_timing[2][192+14].t_rxd2[1][2] = 2332ns;
slave_timing[2][192+14].t_rxd2[2][1] = 2064ns;

slave_timing[2][192+15].info_corner          = 3;
slave_timing[2][192+15].info_temp__j__       = -40;
slave_timing[2][192+15].info_i__quite_rec__  = 0.003000000;
slave_timing[2][192+15].info_dtr__ib__       = 1;
slave_timing[2][192+15].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+15].info_i__max_slave__  = 0.025000000;
slave_timing[2][192+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][192+15].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+15].t_rxd1[0][1] = 2223ns;
slave_timing[2][192+15].t_rxd1[1][0] = 2311ns;
slave_timing[2][192+15].t_rxd1[0][2] = 1698ns;
slave_timing[2][192+15].t_rxd1[2][0] = 2776ns;
slave_timing[2][192+15].t_rxd2[0][2] = 2604ns;
slave_timing[2][192+15].t_rxd2[2][0] = 1726ns;
slave_timing[2][192+15].t_rxd2[1][2] = 2123ns;
slave_timing[2][192+15].t_rxd2[2][1] = 2269ns;

slave_timing[2][192+16].info_corner          = 3;
slave_timing[2][192+16].info_temp__j__       = -40;
slave_timing[2][192+16].info_i__quite_rec__  = 0.000000000;
slave_timing[2][192+16].info_dtr__ib__       = -1;
slave_timing[2][192+16].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+16].info_i__max_slave__  = 0.023000000;
slave_timing[2][192+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][192+16].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+16].t_rxd1[0][1] = 2193ns;
slave_timing[2][192+16].t_rxd1[1][0] = 2205ns;
slave_timing[2][192+16].t_rxd1[0][2] = 1657ns;
slave_timing[2][192+16].t_rxd1[2][0] = 2679ns;
slave_timing[2][192+16].t_rxd2[0][2] = 2644ns;
slave_timing[2][192+16].t_rxd2[2][0] = 1671ns;
slave_timing[2][192+16].t_rxd2[1][2] = 2165ns;
slave_timing[2][192+16].t_rxd2[2][1] = 2210ns;

slave_timing[2][192+17].info_corner          = 3;
slave_timing[2][192+17].info_temp__j__       = -40;
slave_timing[2][192+17].info_i__quite_rec__  = 0.000000000;
slave_timing[2][192+17].info_dtr__ib__       = -1;
slave_timing[2][192+17].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+17].info_i__max_slave__  = 0.025000000;
slave_timing[2][192+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][192+17].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+17].t_rxd1[0][1] = 2108ns;
slave_timing[2][192+17].t_rxd1[1][0] = 2269ns;
slave_timing[2][192+17].t_rxd1[0][2] = 1590ns;
slave_timing[2][192+17].t_rxd1[2][0] = 2733ns;
slave_timing[2][192+17].t_rxd2[0][2] = 2479ns;
slave_timing[2][192+17].t_rxd2[2][0] = 1784ns;
slave_timing[2][192+17].t_rxd2[1][2] = 1936ns;
slave_timing[2][192+17].t_rxd2[2][1] = 2432ns;

slave_timing[2][192+18].info_corner          = 3;
slave_timing[2][192+18].info_temp__j__       = -40;
slave_timing[2][192+18].info_i__quite_rec__  = 0.000000000;
slave_timing[2][192+18].info_dtr__ib__       = 1;
slave_timing[2][192+18].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+18].info_i__max_slave__  = 0.023000000;
slave_timing[2][192+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][192+18].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+18].t_rxd1[0][1] = 2252ns;
slave_timing[2][192+18].t_rxd1[1][0] = 2148ns;
slave_timing[2][192+18].t_rxd1[0][2] = 1690ns;
slave_timing[2][192+18].t_rxd1[2][0] = 2645ns;
slave_timing[2][192+18].t_rxd2[0][2] = 2776ns;
slave_timing[2][192+18].t_rxd2[2][0] = 1551ns;
slave_timing[2][192+18].t_rxd2[1][2] = 2359ns;
slave_timing[2][192+18].t_rxd2[2][1] = 2024ns;

slave_timing[2][192+19].info_corner          = 3;
slave_timing[2][192+19].info_temp__j__       = -40;
slave_timing[2][192+19].info_i__quite_rec__  = 0.000000000;
slave_timing[2][192+19].info_dtr__ib__       = 1;
slave_timing[2][192+19].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+19].info_i__max_slave__  = 0.025000000;
slave_timing[2][192+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][192+19].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+19].t_rxd1[0][1] = 2180ns;
slave_timing[2][192+19].t_rxd1[1][0] = 2214ns;
slave_timing[2][192+19].t_rxd1[0][2] = 1645ns;
slave_timing[2][192+19].t_rxd1[2][0] = 2697ns;
slave_timing[2][192+19].t_rxd2[0][2] = 2602ns;
slave_timing[2][192+19].t_rxd2[2][0] = 1698ns;
slave_timing[2][192+19].t_rxd2[1][2] = 2078ns;
slave_timing[2][192+19].t_rxd2[2][1] = 2254ns;

slave_timing[2][192+20].info_corner          = 3;
slave_timing[2][192+20].info_temp__j__       = -40;
slave_timing[2][192+20].info_i__quite_rec__  = 0.000000000;
slave_timing[2][192+20].info_dtr__ib__       = -1;
slave_timing[2][192+20].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+20].info_i__max_slave__  = 0.023000000;
slave_timing[2][192+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][192+20].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+20].t_rxd1[0][1] = 2278ns;
slave_timing[2][192+20].t_rxd1[1][0] = 2275ns;
slave_timing[2][192+20].t_rxd1[0][2] = 1731ns;
slave_timing[2][192+20].t_rxd1[2][0] = 2759ns;
slave_timing[2][192+20].t_rxd2[0][2] = 2653ns;
slave_timing[2][192+20].t_rxd2[2][0] = 1683ns;
slave_timing[2][192+20].t_rxd2[1][2] = 2171ns;
slave_timing[2][192+20].t_rxd2[2][1] = 2215ns;

slave_timing[2][192+21].info_corner          = 3;
slave_timing[2][192+21].info_temp__j__       = -40;
slave_timing[2][192+21].info_i__quite_rec__  = 0.000000000;
slave_timing[2][192+21].info_dtr__ib__       = -1;
slave_timing[2][192+21].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+21].info_i__max_slave__  = 0.025000000;
slave_timing[2][192+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][192+21].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+21].t_rxd1[0][1] = 2200ns;
slave_timing[2][192+21].t_rxd1[1][0] = 2349ns;
slave_timing[2][192+21].t_rxd1[0][2] = 1685ns;
slave_timing[2][192+21].t_rxd1[2][0] = 2802ns;
slave_timing[2][192+21].t_rxd2[0][2] = 2513ns;
slave_timing[2][192+21].t_rxd2[2][0] = 1798ns;
slave_timing[2][192+21].t_rxd2[1][2] = 1946ns;
slave_timing[2][192+21].t_rxd2[2][1] = 2421ns;

slave_timing[2][192+22].info_corner          = 3;
slave_timing[2][192+22].info_temp__j__       = -40;
slave_timing[2][192+22].info_i__quite_rec__  = 0.000000000;
slave_timing[2][192+22].info_dtr__ib__       = 1;
slave_timing[2][192+22].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+22].info_i__max_slave__  = 0.023000000;
slave_timing[2][192+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][192+22].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+22].t_rxd1[0][1] = 2334ns;
slave_timing[2][192+22].t_rxd1[1][0] = 2223ns;
slave_timing[2][192+22].t_rxd1[0][2] = 1762ns;
slave_timing[2][192+22].t_rxd1[2][0] = 2713ns;
slave_timing[2][192+22].t_rxd2[0][2] = 2784ns;
slave_timing[2][192+22].t_rxd2[2][0] = 1569ns;
slave_timing[2][192+22].t_rxd2[1][2] = 2363ns;
slave_timing[2][192+22].t_rxd2[2][1] = 1999ns;

slave_timing[2][192+23].info_corner          = 3;
slave_timing[2][192+23].info_temp__j__       = -40;
slave_timing[2][192+23].info_i__quite_rec__  = 0.000000000;
slave_timing[2][192+23].info_dtr__ib__       = 1;
slave_timing[2][192+23].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+23].info_i__max_slave__  = 0.025000000;
slave_timing[2][192+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][192+23].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+23].t_rxd1[0][1] = 2232ns;
slave_timing[2][192+23].t_rxd1[1][0] = 2290ns;
slave_timing[2][192+23].t_rxd1[0][2] = 1707ns;
slave_timing[2][192+23].t_rxd1[2][0] = 2762ns;
slave_timing[2][192+23].t_rxd2[0][2] = 2616ns;
slave_timing[2][192+23].t_rxd2[2][0] = 1710ns;
slave_timing[2][192+23].t_rxd2[1][2] = 2111ns;
slave_timing[2][192+23].t_rxd2[2][1] = 2269ns;

slave_timing[2][192+24].info_corner          = 3;
slave_timing[2][192+24].info_temp__j__       = -40;
slave_timing[2][192+24].info_i__quite_rec__  = 0.040000000;
slave_timing[2][192+24].info_dtr__ib__       = -1;
slave_timing[2][192+24].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+24].info_i__max_slave__  = 0.023000000;
slave_timing[2][192+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][192+24].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+24].t_rxd1[0][1] = 2193ns;
slave_timing[2][192+24].t_rxd1[1][0] = 2179ns;
slave_timing[2][192+24].t_rxd1[0][2] = 1652ns;
slave_timing[2][192+24].t_rxd1[2][0] = 2668ns;
slave_timing[2][192+24].t_rxd2[0][2] = 2648ns;
slave_timing[2][192+24].t_rxd2[2][0] = 1661ns;
slave_timing[2][192+24].t_rxd2[1][2] = 2163ns;
slave_timing[2][192+24].t_rxd2[2][1] = 2197ns;

slave_timing[2][192+25].info_corner          = 3;
slave_timing[2][192+25].info_temp__j__       = -40;
slave_timing[2][192+25].info_i__quite_rec__  = 0.040000000;
slave_timing[2][192+25].info_dtr__ib__       = -1;
slave_timing[2][192+25].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+25].info_i__max_slave__  = 0.025000000;
slave_timing[2][192+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][192+25].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+25].t_rxd1[0][1] = 2107ns;
slave_timing[2][192+25].t_rxd1[1][0] = 2245ns;
slave_timing[2][192+25].t_rxd1[0][2] = 1600ns;
slave_timing[2][192+25].t_rxd1[2][0] = 2718ns;
slave_timing[2][192+25].t_rxd2[0][2] = 2497ns;
slave_timing[2][192+25].t_rxd2[2][0] = 1778ns;
slave_timing[2][192+25].t_rxd2[1][2] = 1941ns;
slave_timing[2][192+25].t_rxd2[2][1] = 2433ns;

slave_timing[2][192+26].info_corner          = 3;
slave_timing[2][192+26].info_temp__j__       = -40;
slave_timing[2][192+26].info_i__quite_rec__  = 0.040000000;
slave_timing[2][192+26].info_dtr__ib__       = 1;
slave_timing[2][192+26].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+26].info_i__max_slave__  = 0.023000000;
slave_timing[2][192+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][192+26].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+26].t_rxd1[0][1] = 2253ns;
slave_timing[2][192+26].t_rxd1[1][0] = 2129ns;
slave_timing[2][192+26].t_rxd1[0][2] = 1659ns;
slave_timing[2][192+26].t_rxd1[2][0] = 2634ns;
slave_timing[2][192+26].t_rxd2[0][2] = 2769ns;
slave_timing[2][192+26].t_rxd2[2][0] = 1561ns;
slave_timing[2][192+26].t_rxd2[1][2] = 2358ns;
slave_timing[2][192+26].t_rxd2[2][1] = 2019ns;

slave_timing[2][192+27].info_corner          = 3;
slave_timing[2][192+27].info_temp__j__       = -40;
slave_timing[2][192+27].info_i__quite_rec__  = 0.040000000;
slave_timing[2][192+27].info_dtr__ib__       = 1;
slave_timing[2][192+27].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+27].info_i__max_slave__  = 0.025000000;
slave_timing[2][192+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][192+27].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+27].t_rxd1[0][1] = 2160ns;
slave_timing[2][192+27].t_rxd1[1][0] = 2204ns;
slave_timing[2][192+27].t_rxd1[0][2] = 1620ns;
slave_timing[2][192+27].t_rxd1[2][0] = 2688ns;
slave_timing[2][192+27].t_rxd2[0][2] = 2582ns;
slave_timing[2][192+27].t_rxd2[2][0] = 1700ns;
slave_timing[2][192+27].t_rxd2[1][2] = 2095ns;
slave_timing[2][192+27].t_rxd2[2][1] = 2265ns;

slave_timing[2][192+28].info_corner          = 3;
slave_timing[2][192+28].info_temp__j__       = -40;
slave_timing[2][192+28].info_i__quite_rec__  = 0.040000000;
slave_timing[2][192+28].info_dtr__ib__       = -1;
slave_timing[2][192+28].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+28].info_i__max_slave__  = 0.023000000;
slave_timing[2][192+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][192+28].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+28].t_rxd1[0][1] = 2240ns;
slave_timing[2][192+28].t_rxd1[1][0] = 2230ns;
slave_timing[2][192+28].t_rxd1[0][2] = 1692ns;
slave_timing[2][192+28].t_rxd1[2][0] = 2714ns;
slave_timing[2][192+28].t_rxd2[0][2] = 2660ns;
slave_timing[2][192+28].t_rxd2[2][0] = 1672ns;
slave_timing[2][192+28].t_rxd2[1][2] = 2179ns;
slave_timing[2][192+28].t_rxd2[2][1] = 2207ns;

slave_timing[2][192+29].info_corner          = 3;
slave_timing[2][192+29].info_temp__j__       = -40;
slave_timing[2][192+29].info_i__quite_rec__  = 0.040000000;
slave_timing[2][192+29].info_dtr__ib__       = -1;
slave_timing[2][192+29].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+29].info_i__max_slave__  = 0.025000000;
slave_timing[2][192+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][192+29].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+29].t_rxd1[0][1] = 2156ns;
slave_timing[2][192+29].t_rxd1[1][0] = 2302ns;
slave_timing[2][192+29].t_rxd1[0][2] = 1644ns;
slave_timing[2][192+29].t_rxd1[2][0] = 2759ns;
slave_timing[2][192+29].t_rxd2[0][2] = 2513ns;
slave_timing[2][192+29].t_rxd2[2][0] = 1795ns;
slave_timing[2][192+29].t_rxd2[1][2] = 1955ns;
slave_timing[2][192+29].t_rxd2[2][1] = 2446ns;

slave_timing[2][192+30].info_corner          = 3;
slave_timing[2][192+30].info_temp__j__       = -40;
slave_timing[2][192+30].info_i__quite_rec__  = 0.040000000;
slave_timing[2][192+30].info_dtr__ib__       = 1;
slave_timing[2][192+30].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+30].info_i__max_slave__  = 0.023000000;
slave_timing[2][192+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][192+30].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+30].t_rxd1[0][1] = 2278ns;
slave_timing[2][192+30].t_rxd1[1][0] = 2179ns;
slave_timing[2][192+30].t_rxd1[0][2] = 1718ns;
slave_timing[2][192+30].t_rxd1[2][0] = 2676ns;
slave_timing[2][192+30].t_rxd2[0][2] = 2782ns;
slave_timing[2][192+30].t_rxd2[2][0] = 1567ns;
slave_timing[2][192+30].t_rxd2[1][2] = 2373ns;
slave_timing[2][192+30].t_rxd2[2][1] = 2043ns;

slave_timing[2][192+31].info_corner          = 3;
slave_timing[2][192+31].info_temp__j__       = -40;
slave_timing[2][192+31].info_i__quite_rec__  = 0.040000000;
slave_timing[2][192+31].info_dtr__ib__       = 1;
slave_timing[2][192+31].info_i__offset_rec__ = 0.000000000;
slave_timing[2][192+31].info_i__max_slave__  = 0.025000000;
slave_timing[2][192+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][192+31].info_r__dsi_bus__    = 5.000;

slave_timing[2][192+31].t_rxd1[0][1] = 2196ns;
slave_timing[2][192+31].t_rxd1[1][0] = 2255ns;
slave_timing[2][192+31].t_rxd1[0][2] = 1674ns;
slave_timing[2][192+31].t_rxd1[2][0] = 2725ns;
slave_timing[2][192+31].t_rxd2[0][2] = 2616ns;
slave_timing[2][192+31].t_rxd2[2][0] = 1713ns;
slave_timing[2][192+31].t_rxd2[1][2] = 2112ns;
slave_timing[2][192+31].t_rxd2[2][1] = 2251ns;

//-----------------------------------------------------------------------------
// Copyright (c) 2023 Elmos SE
// Author     : Eugene - Easy UVM Generator
//
// Description: This file has been generated automatically by Eugene
//				This file should not be modified manually. 
//-----------------------------------------------------------------------------
`ifndef ELIP_BUS_MONITOR_SV
`define ELIP_BUS_MONITOR_SV

class elip_bus_monitor extends uvm_monitor;

	`uvm_component_utils(elip_bus_monitor)
	
	virtual	elip_bus_if vif;

  	elip_bus_config m_config;

  	uvm_analysis_port #(elip_tr) analysis_port;

  	elip_tr m_trans;

  	function new(string name, uvm_component parent);
  		super.new(name, parent);
  		analysis_port = new("analysis_port", this);
	endfunction
		
	// Methods run_phase, and do_mon generated by setting monitor_inc in file spi.tpl
	task run_phase(uvm_phase phase);
		`uvm_info(get_type_name(), "run_phase", UVM_HIGH)
		m_trans = elip_tr::type_id::create("m_trans");
		do_mon();
	endtask
	
	`include "includes/elip_monitor_inc.sv"
	
	// You can insert code here by setting monitor_inc_inside_class in file elip_bus.tpl
	
endclass

// You can insert code here by setting monitor_inc_after_class in file elip_bus.tpl

`endif

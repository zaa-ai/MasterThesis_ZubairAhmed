
slave_timing[1][32+0].info_corner          = 2;
slave_timing[1][32+0].info_temp__j__       = 125;
slave_timing[1][32+0].info_i__quite_rec__  = 0.006000000;
slave_timing[1][32+0].info_dtr__ib__       = -1;
slave_timing[1][32+0].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+0].info_i__max_slave__  = 0.023000000;
slave_timing[1][32+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][32+0].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+0].t_rxd1[0][1] = 1671ns;
slave_timing[1][32+0].t_rxd1[1][0] = 1689ns;
slave_timing[1][32+0].t_rxd1[0][2] = 1262ns;
slave_timing[1][32+0].t_rxd1[2][0] = 2029ns;
slave_timing[1][32+0].t_rxd2[0][2] = 1998ns;
slave_timing[1][32+0].t_rxd2[2][0] = 1268ns;
slave_timing[1][32+0].t_rxd2[1][2] = 1661ns;
slave_timing[1][32+0].t_rxd2[2][1] = 1669ns;

slave_timing[1][32+1].info_corner          = 2;
slave_timing[1][32+1].info_temp__j__       = 125;
slave_timing[1][32+1].info_i__quite_rec__  = 0.006000000;
slave_timing[1][32+1].info_dtr__ib__       = -1;
slave_timing[1][32+1].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+1].info_i__max_slave__  = 0.025000000;
slave_timing[1][32+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][32+1].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+1].t_rxd1[0][1] = 1610ns;
slave_timing[1][32+1].t_rxd1[1][0] = 1736ns;
slave_timing[1][32+1].t_rxd1[0][2] = 1226ns;
slave_timing[1][32+1].t_rxd1[2][0] = 2061ns;
slave_timing[1][32+1].t_rxd2[0][2] = 1880ns;
slave_timing[1][32+1].t_rxd2[2][0] = 1348ns;
slave_timing[1][32+1].t_rxd2[1][2] = 1488ns;
slave_timing[1][32+1].t_rxd2[2][1] = 1838ns;

slave_timing[1][32+2].info_corner          = 2;
slave_timing[1][32+2].info_temp__j__       = 125;
slave_timing[1][32+2].info_i__quite_rec__  = 0.006000000;
slave_timing[1][32+2].info_dtr__ib__       = 1;
slave_timing[1][32+2].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+2].info_i__max_slave__  = 0.023000000;
slave_timing[1][32+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][32+2].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+2].t_rxd1[0][1] = 1703ns;
slave_timing[1][32+2].t_rxd1[1][0] = 1647ns;
slave_timing[1][32+2].t_rxd1[0][2] = 1274ns;
slave_timing[1][32+2].t_rxd1[2][0] = 1991ns;
slave_timing[1][32+2].t_rxd2[0][2] = 2098ns;
slave_timing[1][32+2].t_rxd2[2][0] = 1193ns;
slave_timing[1][32+2].t_rxd2[1][2] = 1806ns;
slave_timing[1][32+2].t_rxd2[2][1] = 1534ns;

slave_timing[1][32+3].info_corner          = 2;
slave_timing[1][32+3].info_temp__j__       = 125;
slave_timing[1][32+3].info_i__quite_rec__  = 0.006000000;
slave_timing[1][32+3].info_dtr__ib__       = 1;
slave_timing[1][32+3].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+3].info_i__max_slave__  = 0.025000000;
slave_timing[1][32+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][32+3].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+3].t_rxd1[0][1] = 1636ns;
slave_timing[1][32+3].t_rxd1[1][0] = 1693ns;
slave_timing[1][32+3].t_rxd1[0][2] = 1239ns;
slave_timing[1][32+3].t_rxd1[2][0] = 2024ns;
slave_timing[1][32+3].t_rxd2[0][2] = 1954ns;
slave_timing[1][32+3].t_rxd2[2][0] = 1281ns;
slave_timing[1][32+3].t_rxd2[1][2] = 1609ns;
slave_timing[1][32+3].t_rxd2[2][1] = 1698ns;

slave_timing[1][32+4].info_corner          = 2;
slave_timing[1][32+4].info_temp__j__       = 125;
slave_timing[1][32+4].info_i__quite_rec__  = 0.006000000;
slave_timing[1][32+4].info_dtr__ib__       = -1;
slave_timing[1][32+4].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+4].info_i__max_slave__  = 0.023000000;
slave_timing[1][32+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][32+4].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+4].t_rxd1[0][1] = 1841ns;
slave_timing[1][32+4].t_rxd1[1][0] = 1819ns;
slave_timing[1][32+4].t_rxd1[0][2] = 1398ns;
slave_timing[1][32+4].t_rxd1[2][0] = 2155ns;
slave_timing[1][32+4].t_rxd2[0][2] = 2035ns;
slave_timing[1][32+4].t_rxd2[2][0] = 1300ns;
slave_timing[1][32+4].t_rxd2[1][2] = 1683ns;
slave_timing[1][32+4].t_rxd2[2][1] = 1693ns;

slave_timing[1][32+5].info_corner          = 2;
slave_timing[1][32+5].info_temp__j__       = 125;
slave_timing[1][32+5].info_i__quite_rec__  = 0.006000000;
slave_timing[1][32+5].info_dtr__ib__       = -1;
slave_timing[1][32+5].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+5].info_i__max_slave__  = 0.025000000;
slave_timing[1][32+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][32+5].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+5].t_rxd1[0][1] = 1771ns;
slave_timing[1][32+5].t_rxd1[1][0] = 1866ns;
slave_timing[1][32+5].t_rxd1[0][2] = 1360ns;
slave_timing[1][32+5].t_rxd1[2][0] = 2184ns;
slave_timing[1][32+5].t_rxd2[0][2] = 1919ns;
slave_timing[1][32+5].t_rxd2[2][0] = 1378ns;
slave_timing[1][32+5].t_rxd2[1][2] = 1535ns;
slave_timing[1][32+5].t_rxd2[2][1] = 1833ns;

slave_timing[1][32+6].info_corner          = 2;
slave_timing[1][32+6].info_temp__j__       = 125;
slave_timing[1][32+6].info_i__quite_rec__  = 0.006000000;
slave_timing[1][32+6].info_dtr__ib__       = 1;
slave_timing[1][32+6].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+6].info_i__max_slave__  = 0.023000000;
slave_timing[1][32+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][32+6].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+6].t_rxd1[0][1] = 1875ns;
slave_timing[1][32+6].t_rxd1[1][0] = 1775ns;
slave_timing[1][32+6].t_rxd1[0][2] = 1412ns;
slave_timing[1][32+6].t_rxd1[2][0] = 2114ns;
slave_timing[1][32+6].t_rxd2[0][2] = 2130ns;
slave_timing[1][32+6].t_rxd2[2][0] = 1220ns;
slave_timing[1][32+6].t_rxd2[1][2] = 1824ns;
slave_timing[1][32+6].t_rxd2[2][1] = 1557ns;

slave_timing[1][32+7].info_corner          = 2;
slave_timing[1][32+7].info_temp__j__       = 125;
slave_timing[1][32+7].info_i__quite_rec__  = 0.006000000;
slave_timing[1][32+7].info_dtr__ib__       = 1;
slave_timing[1][32+7].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+7].info_i__max_slave__  = 0.025000000;
slave_timing[1][32+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][32+7].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+7].t_rxd1[0][1] = 1802ns;
slave_timing[1][32+7].t_rxd1[1][0] = 1824ns;
slave_timing[1][32+7].t_rxd1[0][2] = 1373ns;
slave_timing[1][32+7].t_rxd1[2][0] = 2147ns;
slave_timing[1][32+7].t_rxd2[0][2] = 1989ns;
slave_timing[1][32+7].t_rxd2[2][0] = 1311ns;
slave_timing[1][32+7].t_rxd2[1][2] = 1629ns;
slave_timing[1][32+7].t_rxd2[2][1] = 1719ns;

slave_timing[1][32+8].info_corner          = 2;
slave_timing[1][32+8].info_temp__j__       = 125;
slave_timing[1][32+8].info_i__quite_rec__  = 0.003000000;
slave_timing[1][32+8].info_dtr__ib__       = -1;
slave_timing[1][32+8].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+8].info_i__max_slave__  = 0.023000000;
slave_timing[1][32+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][32+8].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+8].t_rxd1[0][1] = 1658ns;
slave_timing[1][32+8].t_rxd1[1][0] = 1665ns;
slave_timing[1][32+8].t_rxd1[0][2] = 1249ns;
slave_timing[1][32+8].t_rxd1[2][0] = 2001ns;
slave_timing[1][32+8].t_rxd2[0][2] = 1988ns;
slave_timing[1][32+8].t_rxd2[2][0] = 1254ns;
slave_timing[1][32+8].t_rxd2[1][2] = 1664ns;
slave_timing[1][32+8].t_rxd2[2][1] = 1645ns;

slave_timing[1][32+9].info_corner          = 2;
slave_timing[1][32+9].info_temp__j__       = 125;
slave_timing[1][32+9].info_i__quite_rec__  = 0.003000000;
slave_timing[1][32+9].info_dtr__ib__       = -1;
slave_timing[1][32+9].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+9].info_i__max_slave__  = 0.025000000;
slave_timing[1][32+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][32+9].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+9].t_rxd1[0][1] = 1592ns;
slave_timing[1][32+9].t_rxd1[1][0] = 1710ns;
slave_timing[1][32+9].t_rxd1[0][2] = 1216ns;
slave_timing[1][32+9].t_rxd1[2][0] = 2032ns;
slave_timing[1][32+9].t_rxd2[0][2] = 1870ns;
slave_timing[1][32+9].t_rxd2[2][0] = 1332ns;
slave_timing[1][32+9].t_rxd2[1][2] = 1492ns;
slave_timing[1][32+9].t_rxd2[2][1] = 1810ns;

slave_timing[1][32+10].info_corner          = 2;
slave_timing[1][32+10].info_temp__j__       = 125;
slave_timing[1][32+10].info_i__quite_rec__  = 0.003000000;
slave_timing[1][32+10].info_dtr__ib__       = 1;
slave_timing[1][32+10].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+10].info_i__max_slave__  = 0.023000000;
slave_timing[1][32+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][32+10].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+10].t_rxd1[0][1] = 1683ns;
slave_timing[1][32+10].t_rxd1[1][0] = 1602ns;
slave_timing[1][32+10].t_rxd1[0][2] = 1256ns;
slave_timing[1][32+10].t_rxd1[2][0] = 1946ns;
slave_timing[1][32+10].t_rxd2[0][2] = 2083ns;
slave_timing[1][32+10].t_rxd2[2][0] = 1177ns;
slave_timing[1][32+10].t_rxd2[1][2] = 1803ns;
slave_timing[1][32+10].t_rxd2[2][1] = 1513ns;

slave_timing[1][32+11].info_corner          = 2;
slave_timing[1][32+11].info_temp__j__       = 125;
slave_timing[1][32+11].info_i__quite_rec__  = 0.003000000;
slave_timing[1][32+11].info_dtr__ib__       = 1;
slave_timing[1][32+11].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+11].info_i__max_slave__  = 0.025000000;
slave_timing[1][32+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][32+11].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+11].t_rxd1[0][1] = 1615ns;
slave_timing[1][32+11].t_rxd1[1][0] = 1648ns;
slave_timing[1][32+11].t_rxd1[0][2] = 1221ns;
slave_timing[1][32+11].t_rxd1[2][0] = 1979ns;
slave_timing[1][32+11].t_rxd2[0][2] = 1938ns;
slave_timing[1][32+11].t_rxd2[2][0] = 1267ns;
slave_timing[1][32+11].t_rxd2[1][2] = 1606ns;
slave_timing[1][32+11].t_rxd2[2][1] = 1678ns;

slave_timing[1][32+12].info_corner          = 2;
slave_timing[1][32+12].info_temp__j__       = 125;
slave_timing[1][32+12].info_i__quite_rec__  = 0.003000000;
slave_timing[1][32+12].info_dtr__ib__       = -1;
slave_timing[1][32+12].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+12].info_i__max_slave__  = 0.023000000;
slave_timing[1][32+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][32+12].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+12].t_rxd1[0][1] = 1839ns;
slave_timing[1][32+12].t_rxd1[1][0] = 1798ns;
slave_timing[1][32+12].t_rxd1[0][2] = 1397ns;
slave_timing[1][32+12].t_rxd1[2][0] = 2125ns;
slave_timing[1][32+12].t_rxd2[0][2] = 2023ns;
slave_timing[1][32+12].t_rxd2[2][0] = 1283ns;
slave_timing[1][32+12].t_rxd2[1][2] = 1684ns;
slave_timing[1][32+12].t_rxd2[2][1] = 1642ns;

slave_timing[1][32+13].info_corner          = 2;
slave_timing[1][32+13].info_temp__j__       = 125;
slave_timing[1][32+13].info_i__quite_rec__  = 0.003000000;
slave_timing[1][32+13].info_dtr__ib__       = -1;
slave_timing[1][32+13].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+13].info_i__max_slave__  = 0.025000000;
slave_timing[1][32+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][32+13].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+13].t_rxd1[0][1] = 1770ns;
slave_timing[1][32+13].t_rxd1[1][0] = 1842ns;
slave_timing[1][32+13].t_rxd1[0][2] = 1343ns;
slave_timing[1][32+13].t_rxd1[2][0] = 2155ns;
slave_timing[1][32+13].t_rxd2[0][2] = 1890ns;
slave_timing[1][32+13].t_rxd2[2][0] = 1362ns;
slave_timing[1][32+13].t_rxd2[1][2] = 1515ns;
slave_timing[1][32+13].t_rxd2[2][1] = 1830ns;

slave_timing[1][32+14].info_corner          = 2;
slave_timing[1][32+14].info_temp__j__       = 125;
slave_timing[1][32+14].info_i__quite_rec__  = 0.003000000;
slave_timing[1][32+14].info_dtr__ib__       = 1;
slave_timing[1][32+14].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+14].info_i__max_slave__  = 0.023000000;
slave_timing[1][32+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][32+14].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+14].t_rxd1[0][1] = 1867ns;
slave_timing[1][32+14].t_rxd1[1][0] = 1733ns;
slave_timing[1][32+14].t_rxd1[0][2] = 1406ns;
slave_timing[1][32+14].t_rxd1[2][0] = 2067ns;
slave_timing[1][32+14].t_rxd2[0][2] = 2111ns;
slave_timing[1][32+14].t_rxd2[2][0] = 1204ns;
slave_timing[1][32+14].t_rxd2[1][2] = 1818ns;
slave_timing[1][32+14].t_rxd2[2][1] = 1537ns;

slave_timing[1][32+15].info_corner          = 2;
slave_timing[1][32+15].info_temp__j__       = 125;
slave_timing[1][32+15].info_i__quite_rec__  = 0.003000000;
slave_timing[1][32+15].info_dtr__ib__       = 1;
slave_timing[1][32+15].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+15].info_i__max_slave__  = 0.025000000;
slave_timing[1][32+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][32+15].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+15].t_rxd1[0][1] = 1792ns;
slave_timing[1][32+15].t_rxd1[1][0] = 1781ns;
slave_timing[1][32+15].t_rxd1[0][2] = 1366ns;
slave_timing[1][32+15].t_rxd1[2][0] = 2100ns;
slave_timing[1][32+15].t_rxd2[0][2] = 1970ns;
slave_timing[1][32+15].t_rxd2[2][0] = 1295ns;
slave_timing[1][32+15].t_rxd2[1][2] = 1628ns;
slave_timing[1][32+15].t_rxd2[2][1] = 1698ns;

slave_timing[1][32+16].info_corner          = 2;
slave_timing[1][32+16].info_temp__j__       = 125;
slave_timing[1][32+16].info_i__quite_rec__  = 0.000000000;
slave_timing[1][32+16].info_dtr__ib__       = -1;
slave_timing[1][32+16].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+16].info_i__max_slave__  = 0.023000000;
slave_timing[1][32+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][32+16].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+16].t_rxd1[0][1] = 1633ns;
slave_timing[1][32+16].t_rxd1[1][0] = 1628ns;
slave_timing[1][32+16].t_rxd1[0][2] = 1230ns;
slave_timing[1][32+16].t_rxd1[2][0] = 1956ns;
slave_timing[1][32+16].t_rxd2[0][2] = 1965ns;
slave_timing[1][32+16].t_rxd2[2][0] = 1238ns;
slave_timing[1][32+16].t_rxd2[1][2] = 1653ns;
slave_timing[1][32+16].t_rxd2[2][1] = 1623ns;

slave_timing[1][32+17].info_corner          = 2;
slave_timing[1][32+17].info_temp__j__       = 125;
slave_timing[1][32+17].info_i__quite_rec__  = 0.000000000;
slave_timing[1][32+17].info_dtr__ib__       = -1;
slave_timing[1][32+17].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+17].info_i__max_slave__  = 0.025000000;
slave_timing[1][32+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][32+17].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+17].t_rxd1[0][1] = 1570ns;
slave_timing[1][32+17].t_rxd1[1][0] = 1670ns;
slave_timing[1][32+17].t_rxd1[0][2] = 1196ns;
slave_timing[1][32+17].t_rxd1[2][0] = 1988ns;
slave_timing[1][32+17].t_rxd2[0][2] = 1846ns;
slave_timing[1][32+17].t_rxd2[2][0] = 1318ns;
slave_timing[1][32+17].t_rxd2[1][2] = 1482ns;
slave_timing[1][32+17].t_rxd2[2][1] = 1785ns;

slave_timing[1][32+18].info_corner          = 2;
slave_timing[1][32+18].info_temp__j__       = 125;
slave_timing[1][32+18].info_i__quite_rec__  = 0.000000000;
slave_timing[1][32+18].info_dtr__ib__       = 1;
slave_timing[1][32+18].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+18].info_i__max_slave__  = 0.023000000;
slave_timing[1][32+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][32+18].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+18].t_rxd1[0][1] = 1660ns;
slave_timing[1][32+18].t_rxd1[1][0] = 1576ns;
slave_timing[1][32+18].t_rxd1[0][2] = 1238ns;
slave_timing[1][32+18].t_rxd1[2][0] = 1908ns;
slave_timing[1][32+18].t_rxd2[0][2] = 2053ns;
slave_timing[1][32+18].t_rxd2[2][0] = 1152ns;
slave_timing[1][32+18].t_rxd2[1][2] = 1781ns;
slave_timing[1][32+18].t_rxd2[2][1] = 1483ns;

slave_timing[1][32+19].info_corner          = 2;
slave_timing[1][32+19].info_temp__j__       = 125;
slave_timing[1][32+19].info_i__quite_rec__  = 0.000000000;
slave_timing[1][32+19].info_dtr__ib__       = 1;
slave_timing[1][32+19].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+19].info_i__max_slave__  = 0.025000000;
slave_timing[1][32+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][32+19].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+19].t_rxd1[0][1] = 1588ns;
slave_timing[1][32+19].t_rxd1[1][0] = 1624ns;
slave_timing[1][32+19].t_rxd1[0][2] = 1202ns;
slave_timing[1][32+19].t_rxd1[2][0] = 1941ns;
slave_timing[1][32+19].t_rxd2[0][2] = 1909ns;
slave_timing[1][32+19].t_rxd2[2][0] = 1245ns;
slave_timing[1][32+19].t_rxd2[1][2] = 1592ns;
slave_timing[1][32+19].t_rxd2[2][1] = 1644ns;

slave_timing[1][32+20].info_corner          = 2;
slave_timing[1][32+20].info_temp__j__       = 125;
slave_timing[1][32+20].info_i__quite_rec__  = 0.000000000;
slave_timing[1][32+20].info_dtr__ib__       = -1;
slave_timing[1][32+20].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+20].info_i__max_slave__  = 0.023000000;
slave_timing[1][32+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][32+20].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+20].t_rxd1[0][1] = 1830ns;
slave_timing[1][32+20].t_rxd1[1][0] = 1754ns;
slave_timing[1][32+20].t_rxd1[0][2] = 1390ns;
slave_timing[1][32+20].t_rxd1[2][0] = 2073ns;
slave_timing[1][32+20].t_rxd2[0][2] = 1994ns;
slave_timing[1][32+20].t_rxd2[2][0] = 1266ns;
slave_timing[1][32+20].t_rxd2[1][2] = 1672ns;
slave_timing[1][32+20].t_rxd2[2][1] = 1641ns;

slave_timing[1][32+21].info_corner          = 2;
slave_timing[1][32+21].info_temp__j__       = 125;
slave_timing[1][32+21].info_i__quite_rec__  = 0.000000000;
slave_timing[1][32+21].info_dtr__ib__       = -1;
slave_timing[1][32+21].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+21].info_i__max_slave__  = 0.025000000;
slave_timing[1][32+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][32+21].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+21].t_rxd1[0][1] = 1761ns;
slave_timing[1][32+21].t_rxd1[1][0] = 1797ns;
slave_timing[1][32+21].t_rxd1[0][2] = 1353ns;
slave_timing[1][32+21].t_rxd1[2][0] = 2105ns;
slave_timing[1][32+21].t_rxd2[0][2] = 1880ns;
slave_timing[1][32+21].t_rxd2[2][0] = 1348ns;
slave_timing[1][32+21].t_rxd2[1][2] = 1526ns;
slave_timing[1][32+21].t_rxd2[2][1] = 1783ns;

slave_timing[1][32+22].info_corner          = 2;
slave_timing[1][32+22].info_temp__j__       = 125;
slave_timing[1][32+22].info_i__quite_rec__  = 0.000000000;
slave_timing[1][32+22].info_dtr__ib__       = 1;
slave_timing[1][32+22].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+22].info_i__max_slave__  = 0.023000000;
slave_timing[1][32+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][32+22].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+22].t_rxd1[0][1] = 1860ns;
slave_timing[1][32+22].t_rxd1[1][0] = 1706ns;
slave_timing[1][32+22].t_rxd1[0][2] = 1400ns;
slave_timing[1][32+22].t_rxd1[2][0] = 2026ns;
slave_timing[1][32+22].t_rxd2[0][2] = 2073ns;
slave_timing[1][32+22].t_rxd2[2][0] = 1182ns;
slave_timing[1][32+22].t_rxd2[1][2] = 1830ns;
slave_timing[1][32+22].t_rxd2[2][1] = 1485ns;

slave_timing[1][32+23].info_corner          = 2;
slave_timing[1][32+23].info_temp__j__       = 125;
slave_timing[1][32+23].info_i__quite_rec__  = 0.000000000;
slave_timing[1][32+23].info_dtr__ib__       = 1;
slave_timing[1][32+23].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+23].info_i__max_slave__  = 0.025000000;
slave_timing[1][32+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][32+23].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+23].t_rxd1[0][1] = 1787ns;
slave_timing[1][32+23].t_rxd1[1][0] = 1751ns;
slave_timing[1][32+23].t_rxd1[0][2] = 1363ns;
slave_timing[1][32+23].t_rxd1[2][0] = 2057ns;
slave_timing[1][32+23].t_rxd2[0][2] = 1938ns;
slave_timing[1][32+23].t_rxd2[2][0] = 1272ns;
slave_timing[1][32+23].t_rxd2[1][2] = 1608ns;
slave_timing[1][32+23].t_rxd2[2][1] = 1644ns;

slave_timing[1][32+24].info_corner          = 2;
slave_timing[1][32+24].info_temp__j__       = 125;
slave_timing[1][32+24].info_i__quite_rec__  = 0.040000000;
slave_timing[1][32+24].info_dtr__ib__       = -1;
slave_timing[1][32+24].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+24].info_i__max_slave__  = 0.023000000;
slave_timing[1][32+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][32+24].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+24].t_rxd1[0][1] = 1664ns;
slave_timing[1][32+24].t_rxd1[1][0] = 1693ns;
slave_timing[1][32+24].t_rxd1[0][2] = 1264ns;
slave_timing[1][32+24].t_rxd1[2][0] = 2034ns;
slave_timing[1][32+24].t_rxd2[0][2] = 2176ns;
slave_timing[1][32+24].t_rxd2[2][0] = 1423ns;
slave_timing[1][32+24].t_rxd2[1][2] = 1846ns;
slave_timing[1][32+24].t_rxd2[2][1] = 1860ns;

slave_timing[1][32+25].info_corner          = 2;
slave_timing[1][32+25].info_temp__j__       = 125;
slave_timing[1][32+25].info_i__quite_rec__  = 0.040000000;
slave_timing[1][32+25].info_dtr__ib__       = -1;
slave_timing[1][32+25].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+25].info_i__max_slave__  = 0.025000000;
slave_timing[1][32+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][32+25].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+25].t_rxd1[0][1] = 1601ns;
slave_timing[1][32+25].t_rxd1[1][0] = 1740ns;
slave_timing[1][32+25].t_rxd1[0][2] = 1229ns;
slave_timing[1][32+25].t_rxd1[2][0] = 2069ns;
slave_timing[1][32+25].t_rxd2[0][2] = 2050ns;
slave_timing[1][32+25].t_rxd2[2][0] = 1509ns;
slave_timing[1][32+25].t_rxd2[1][2] = 1671ns;
slave_timing[1][32+25].t_rxd2[2][1] = 2017ns;

slave_timing[1][32+26].info_corner          = 2;
slave_timing[1][32+26].info_temp__j__       = 125;
slave_timing[1][32+26].info_i__quite_rec__  = 0.040000000;
slave_timing[1][32+26].info_dtr__ib__       = 1;
slave_timing[1][32+26].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+26].info_i__max_slave__  = 0.023000000;
slave_timing[1][32+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][32+26].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+26].t_rxd1[0][1] = 1732ns;
slave_timing[1][32+26].t_rxd1[1][0] = 1637ns;
slave_timing[1][32+26].t_rxd1[0][2] = 1296ns;
slave_timing[1][32+26].t_rxd1[2][0] = 1991ns;
slave_timing[1][32+26].t_rxd2[0][2] = 2305ns;
slave_timing[1][32+26].t_rxd2[2][0] = 1336ns;
slave_timing[1][32+26].t_rxd2[1][2] = 2021ns;
slave_timing[1][32+26].t_rxd2[2][1] = 1702ns;

slave_timing[1][32+27].info_corner          = 2;
slave_timing[1][32+27].info_temp__j__       = 125;
slave_timing[1][32+27].info_i__quite_rec__  = 0.040000000;
slave_timing[1][32+27].info_dtr__ib__       = 1;
slave_timing[1][32+27].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+27].info_i__max_slave__  = 0.025000000;
slave_timing[1][32+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][32+27].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+27].t_rxd1[0][1] = 1660ns;
slave_timing[1][32+27].t_rxd1[1][0] = 1688ns;
slave_timing[1][32+27].t_rxd1[0][2] = 1261ns;
slave_timing[1][32+27].t_rxd1[2][0] = 2032ns;
slave_timing[1][32+27].t_rxd2[0][2] = 2150ns;
slave_timing[1][32+27].t_rxd2[2][0] = 1431ns;
slave_timing[1][32+27].t_rxd2[1][2] = 1814ns;
slave_timing[1][32+27].t_rxd2[2][1] = 1883ns;

slave_timing[1][32+28].info_corner          = 2;
slave_timing[1][32+28].info_temp__j__       = 125;
slave_timing[1][32+28].info_i__quite_rec__  = 0.040000000;
slave_timing[1][32+28].info_dtr__ib__       = -1;
slave_timing[1][32+28].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+28].info_i__max_slave__  = 0.023000000;
slave_timing[1][32+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][32+28].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+28].t_rxd1[0][1] = 1736ns;
slave_timing[1][32+28].t_rxd1[1][0] = 1737ns;
slave_timing[1][32+28].t_rxd1[0][2] = 1344ns;
slave_timing[1][32+28].t_rxd1[2][0] = 2405ns;
slave_timing[1][32+28].t_rxd2[0][2] = 2676ns;
slave_timing[1][32+28].t_rxd2[2][0] = 1903ns;
slave_timing[1][32+28].t_rxd2[1][2] = 2399ns;
slave_timing[1][32+28].t_rxd2[2][1] = 2617ns;

slave_timing[1][32+29].info_corner          = 2;
slave_timing[1][32+29].info_temp__j__       = 125;
slave_timing[1][32+29].info_i__quite_rec__  = 0.040000000;
slave_timing[1][32+29].info_dtr__ib__       = -1;
slave_timing[1][32+29].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+29].info_i__max_slave__  = 0.025000000;
slave_timing[1][32+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][32+29].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+29].t_rxd1[0][1] = 1673ns;
slave_timing[1][32+29].t_rxd1[1][0] = 1783ns;
slave_timing[1][32+29].t_rxd1[0][2] = 1312ns;
slave_timing[1][32+29].t_rxd1[2][0] = 2509ns;
slave_timing[1][32+29].t_rxd2[0][2] = 2489ns;
slave_timing[1][32+29].t_rxd2[2][0] = 2038ns;
slave_timing[1][32+29].t_rxd2[1][2] = 2166ns;
slave_timing[1][32+29].t_rxd2[2][1] = 3007ns;

slave_timing[1][32+30].info_corner          = 2;
slave_timing[1][32+30].info_temp__j__       = 125;
slave_timing[1][32+30].info_i__quite_rec__  = 0.040000000;
slave_timing[1][32+30].info_dtr__ib__       = 1;
slave_timing[1][32+30].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+30].info_i__max_slave__  = 0.023000000;
slave_timing[1][32+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][32+30].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+30].t_rxd1[0][1] = 1796ns;
slave_timing[1][32+30].t_rxd1[1][0] = 1683ns;
slave_timing[1][32+30].t_rxd1[0][2] = 1374ns;
slave_timing[1][32+30].t_rxd1[2][0] = 2304ns;
slave_timing[1][32+30].t_rxd2[0][2] = 2889ns;
slave_timing[1][32+30].t_rxd2[2][0] = 1771ns;
slave_timing[1][32+30].t_rxd2[1][2] = 2642ns;
slave_timing[1][32+30].t_rxd2[2][1] = 2330ns;

slave_timing[1][32+31].info_corner          = 2;
slave_timing[1][32+31].info_temp__j__       = 125;
slave_timing[1][32+31].info_i__quite_rec__  = 0.040000000;
slave_timing[1][32+31].info_dtr__ib__       = 1;
slave_timing[1][32+31].info_i__offset_rec__ = 0.000000000;
slave_timing[1][32+31].info_i__max_slave__  = 0.025000000;
slave_timing[1][32+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][32+31].info_r__dsi_bus__    = 5.000;

slave_timing[1][32+31].t_rxd1[0][1] = 1728ns;
slave_timing[1][32+31].t_rxd1[1][0] = 1725ns;
slave_timing[1][32+31].t_rxd1[0][2] = 1337ns;
slave_timing[1][32+31].t_rxd1[2][0] = 2406ns;
slave_timing[1][32+31].t_rxd2[0][2] = 2638ns;
slave_timing[1][32+31].t_rxd2[2][0] = 1917ns;
slave_timing[1][32+31].t_rxd2[1][2] = 2353ns;
slave_timing[1][32+31].t_rxd2[2][1] = 2666ns;

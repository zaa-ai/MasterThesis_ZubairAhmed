// Denso Waveshape reset values
wave_luts[0][0]  <=5'h1f;
wave_luts[0][1]  <=5'h1f;
wave_luts[0][2]  <=5'h1f;
wave_luts[0][3]  <=5'h1f;
wave_luts[0][4]  <=5'h1e;
wave_luts[0][5]  <=5'h1f;
wave_luts[0][6]  <=5'h1e;
wave_luts[0][7]  <=5'h1f;
wave_luts[0][8]  <=5'h1e;
wave_luts[0][9]  <=5'h1e;
wave_luts[0][10] <=5'h1e;
wave_luts[0][11] <=5'h1e;
wave_luts[0][12] <=5'h1d;
wave_luts[0][13] <=5'h1d;
wave_luts[0][14] <=5'h1c;
wave_luts[0][15] <=5'h1c;
wave_luts[0][16] <=5'h1c;
wave_luts[0][17] <=5'h1b;
wave_luts[0][18] <=5'h1a;
wave_luts[0][19] <=5'h1a;
wave_luts[0][20] <=5'h19;
wave_luts[0][21] <=5'h19;
wave_luts[0][22] <=5'h18;
wave_luts[0][23] <=5'h17;
wave_luts[0][24] <=5'h17;
wave_luts[0][25] <=5'h16;
wave_luts[0][26] <=5'h15;
wave_luts[0][27] <=5'h14;
wave_luts[0][28] <=5'h14;
wave_luts[0][29] <=5'h13;
wave_luts[0][30] <=5'h12;
wave_luts[0][31] <=5'h11;
wave_luts[0][32] <=5'h10;
wave_luts[0][33] <=5'h0f;
wave_luts[0][34] <=5'h0e;
wave_luts[0][35] <=5'h0d;
wave_luts[0][36] <=5'h0c;
wave_luts[0][37] <=5'h0b;
wave_luts[0][38] <=5'h0b;
wave_luts[0][39] <=5'h0a;
wave_luts[0][40] <=5'h09;
wave_luts[0][41] <=5'h08;
wave_luts[0][42] <=5'h08;
wave_luts[0][43] <=5'h07;
wave_luts[0][44] <=5'h06;
wave_luts[0][45] <=5'h06;
wave_luts[0][46] <=5'h05;
wave_luts[0][47] <=5'h05;
wave_luts[0][48] <=5'h04;
wave_luts[0][49] <=5'h03;
wave_luts[0][50] <=5'h03;
wave_luts[0][51] <=5'h03;
wave_luts[0][52] <=5'h02;
wave_luts[0][53] <=5'h02;
wave_luts[0][54] <=5'h01;
wave_luts[0][55] <=5'h01;
wave_luts[0][56] <=5'h01;
wave_luts[0][57] <=5'h01;
wave_luts[0][58] <=5'h00;
wave_luts[0][59] <=5'h00;
wave_luts[0][60] <=5'h00;
wave_luts[0][61] <=5'h00;
wave_luts[0][62] <=5'h00;
wave_luts[0][63] <=5'h00;
wave_luts[0][64] <=5'h00;
wave_luts[0][65] <=5'h00;
wave_luts[0][66] <=5'h00;
wave_luts[0][67] <=5'h00;
wave_luts[0][68] <=5'h00;
wave_luts[0][69] <=5'h00;
wave_luts[0][70] <=5'h00;
wave_luts[0][71] <=5'h00;

wave_luts[1][0]  <=5'h00;
wave_luts[1][1]  <=5'h00;
wave_luts[1][2]  <=5'h00;
wave_luts[1][3]  <=5'h00;
wave_luts[1][4]  <=5'h00;
wave_luts[1][5]  <=5'h00;
wave_luts[1][6]  <=5'h00;
wave_luts[1][7]  <=5'h01;
wave_luts[1][8]  <=5'h00;
wave_luts[1][9]  <=5'h01;
wave_luts[1][10] <=5'h01;
wave_luts[1][11] <=5'h02;
wave_luts[1][12] <=5'h01;
wave_luts[1][13] <=5'h02;
wave_luts[1][14] <=5'h02;
wave_luts[1][15] <=5'h03;
wave_luts[1][16] <=5'h03;
wave_luts[1][17] <=5'h04;
wave_luts[1][18] <=5'h04;
wave_luts[1][19] <=5'h05;
wave_luts[1][20] <=5'h05;
wave_luts[1][21] <=5'h06;
wave_luts[1][22] <=5'h06;
wave_luts[1][23] <=5'h07;
wave_luts[1][24] <=5'h08;
wave_luts[1][25] <=5'h08;
wave_luts[1][26] <=5'h09;
wave_luts[1][27] <=5'h0a;
wave_luts[1][28] <=5'h0a;
wave_luts[1][29] <=5'h0b;
wave_luts[1][30] <=5'h0c;
wave_luts[1][31] <=5'h0d;
wave_luts[1][32] <=5'h0e;
wave_luts[1][33] <=5'h0f;
wave_luts[1][34] <=5'h10;
wave_luts[1][35] <=5'h10;
wave_luts[1][36] <=5'h11;
wave_luts[1][37] <=5'h12;
wave_luts[1][38] <=5'h13;
wave_luts[1][39] <=5'h14;
wave_luts[1][40] <=5'h15;
wave_luts[1][41] <=5'h15;
wave_luts[1][42] <=5'h16;
wave_luts[1][43] <=5'h17;
wave_luts[1][44] <=5'h17;
wave_luts[1][45] <=5'h18;
wave_luts[1][46] <=5'h19;
wave_luts[1][47] <=5'h19;
wave_luts[1][48] <=5'h1a;
wave_luts[1][49] <=5'h1a;
wave_luts[1][50] <=5'h1b;
wave_luts[1][51] <=5'h1b;
wave_luts[1][52] <=5'h1c;
wave_luts[1][53] <=5'h1c;
wave_luts[1][54] <=5'h1d;
wave_luts[1][55] <=5'h1d;
wave_luts[1][56] <=5'h1d;
wave_luts[1][57] <=5'h1e;
wave_luts[1][58] <=5'h1e;
wave_luts[1][59] <=5'h1e;
wave_luts[1][60] <=5'h1f;
wave_luts[1][61] <=5'h1f;
wave_luts[1][62] <=5'h1f;
wave_luts[1][63] <=5'h1f;
wave_luts[1][64] <=5'h1f;
wave_luts[1][65] <=5'h1f;
wave_luts[1][66] <=5'h1f;
wave_luts[1][67] <=5'h1f;
wave_luts[1][68] <=5'h1f;
wave_luts[1][69] <=5'h1f;
wave_luts[1][70] <=5'h1f;
wave_luts[1][71] <=5'h1f;

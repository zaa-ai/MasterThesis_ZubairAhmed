/**
 * Package: common_env_pkg
 *
 * Common package for class based items
 */
package common_env_pkg;

endpackage



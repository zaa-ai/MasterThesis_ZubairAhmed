/**
 * Interface: dsi_logic_if
 * 
 * TODO: Add interface documentation
 */
interface dsi_logic_if import project_pkg::*; ();
	
	dsi_logic_t	D;

endinterface

/* ###   interface instances   ###################################################### */

supply_registers_TRIM_IREF_if supply_registers_TRIM_IREF (); 
supply_registers_TRIM_OT_if supply_registers_TRIM_OT (); 
supply_registers_SUP_IRQ_STAT_if supply_registers_SUP_IRQ_STAT (); 
supply_registers_SUP_IRQ_MASK_if supply_registers_SUP_IRQ_MASK (); 
supply_registers_SUP_HW_CTRL_if supply_registers_SUP_HW_CTRL (); 
supply_registers_SUP_STAT_if supply_registers_SUP_STAT (); 
supply_registers_SUP_CTRL_if supply_registers_SUP_CTRL (); 
supply_registers_IO_CTRL_if supply_registers_IO_CTRL (); 



slave_timing[1][224+0].info_corner          = 4;
slave_timing[1][224+0].info_temp__j__       = -40;
slave_timing[1][224+0].info_i__quite_rec__  = 0.006000000;
slave_timing[1][224+0].info_dtr__ib__       = -1;
slave_timing[1][224+0].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+0].info_i__max_slave__  = 0.023000000;
slave_timing[1][224+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][224+0].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+0].t_rxd1[0][1] = 1700ns;
slave_timing[1][224+0].t_rxd1[1][0] = 1680ns;
slave_timing[1][224+0].t_rxd1[0][2] = 1274ns;
slave_timing[1][224+0].t_rxd1[2][0] = 2054ns;
slave_timing[1][224+0].t_rxd2[0][2] = 2059ns;
slave_timing[1][224+0].t_rxd2[2][0] = 1257ns;
slave_timing[1][224+0].t_rxd2[1][2] = 1693ns;
slave_timing[1][224+0].t_rxd2[2][1] = 1662ns;

slave_timing[1][224+1].info_corner          = 4;
slave_timing[1][224+1].info_temp__j__       = -40;
slave_timing[1][224+1].info_i__quite_rec__  = 0.006000000;
slave_timing[1][224+1].info_dtr__ib__       = -1;
slave_timing[1][224+1].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+1].info_i__max_slave__  = 0.025000000;
slave_timing[1][224+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][224+1].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+1].t_rxd1[0][1] = 1636ns;
slave_timing[1][224+1].t_rxd1[1][0] = 1730ns;
slave_timing[1][224+1].t_rxd1[0][2] = 1239ns;
slave_timing[1][224+1].t_rxd1[2][0] = 2089ns;
slave_timing[1][224+1].t_rxd2[0][2] = 1931ns;
slave_timing[1][224+1].t_rxd2[2][0] = 1344ns;
slave_timing[1][224+1].t_rxd2[1][2] = 1511ns;
slave_timing[1][224+1].t_rxd2[2][1] = 1838ns;

slave_timing[1][224+2].info_corner          = 4;
slave_timing[1][224+2].info_temp__j__       = -40;
slave_timing[1][224+2].info_i__quite_rec__  = 0.006000000;
slave_timing[1][224+2].info_dtr__ib__       = 1;
slave_timing[1][224+2].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+2].info_i__max_slave__  = 0.023000000;
slave_timing[1][224+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][224+2].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+2].t_rxd1[0][1] = 1743ns;
slave_timing[1][224+2].t_rxd1[1][0] = 1651ns;
slave_timing[1][224+2].t_rxd1[0][2] = 1297ns;
slave_timing[1][224+2].t_rxd1[2][0] = 2032ns;
slave_timing[1][224+2].t_rxd2[0][2] = 2158ns;
slave_timing[1][224+2].t_rxd2[2][0] = 1196ns;
slave_timing[1][224+2].t_rxd2[1][2] = 1826ns;
slave_timing[1][224+2].t_rxd2[2][1] = 1550ns;

slave_timing[1][224+3].info_corner          = 4;
slave_timing[1][224+3].info_temp__j__       = -40;
slave_timing[1][224+3].info_i__quite_rec__  = 0.006000000;
slave_timing[1][224+3].info_dtr__ib__       = 1;
slave_timing[1][224+3].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+3].info_i__max_slave__  = 0.025000000;
slave_timing[1][224+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][224+3].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+3].t_rxd1[0][1] = 1672ns;
slave_timing[1][224+3].t_rxd1[1][0] = 1703ns;
slave_timing[1][224+3].t_rxd1[0][2] = 1255ns;
slave_timing[1][224+3].t_rxd1[2][0] = 2068ns;
slave_timing[1][224+3].t_rxd2[0][2] = 2005ns;
slave_timing[1][224+3].t_rxd2[2][0] = 1288ns;
slave_timing[1][224+3].t_rxd2[1][2] = 1620ns;
slave_timing[1][224+3].t_rxd2[2][1] = 1705ns;

slave_timing[1][224+4].info_corner          = 4;
slave_timing[1][224+4].info_temp__j__       = -40;
slave_timing[1][224+4].info_i__quite_rec__  = 0.006000000;
slave_timing[1][224+4].info_dtr__ib__       = -1;
slave_timing[1][224+4].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+4].info_i__max_slave__  = 0.023000000;
slave_timing[1][224+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][224+4].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+4].t_rxd1[0][1] = 1781ns;
slave_timing[1][224+4].t_rxd1[1][0] = 1750ns;
slave_timing[1][224+4].t_rxd1[0][2] = 1336ns;
slave_timing[1][224+4].t_rxd1[2][0] = 2120ns;
slave_timing[1][224+4].t_rxd2[0][2] = 2077ns;
slave_timing[1][224+4].t_rxd2[2][0] = 1271ns;
slave_timing[1][224+4].t_rxd2[1][2] = 1704ns;
slave_timing[1][224+4].t_rxd2[2][1] = 1673ns;

slave_timing[1][224+5].info_corner          = 4;
slave_timing[1][224+5].info_temp__j__       = -40;
slave_timing[1][224+5].info_i__quite_rec__  = 0.006000000;
slave_timing[1][224+5].info_dtr__ib__       = -1;
slave_timing[1][224+5].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+5].info_i__max_slave__  = 0.025000000;
slave_timing[1][224+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][224+5].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+5].t_rxd1[0][1] = 1712ns;
slave_timing[1][224+5].t_rxd1[1][0] = 1800ns;
slave_timing[1][224+5].t_rxd1[0][2] = 1299ns;
slave_timing[1][224+5].t_rxd1[2][0] = 2155ns;
slave_timing[1][224+5].t_rxd2[0][2] = 1952ns;
slave_timing[1][224+5].t_rxd2[2][0] = 1357ns;
slave_timing[1][224+5].t_rxd2[1][2] = 1523ns;
slave_timing[1][224+5].t_rxd2[2][1] = 1846ns;

slave_timing[1][224+6].info_corner          = 4;
slave_timing[1][224+6].info_temp__j__       = -40;
slave_timing[1][224+6].info_i__quite_rec__  = 0.006000000;
slave_timing[1][224+6].info_dtr__ib__       = 1;
slave_timing[1][224+6].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+6].info_i__max_slave__  = 0.023000000;
slave_timing[1][224+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][224+6].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+6].t_rxd1[0][1] = 1815ns;
slave_timing[1][224+6].t_rxd1[1][0] = 1714ns;
slave_timing[1][224+6].t_rxd1[0][2] = 1353ns;
slave_timing[1][224+6].t_rxd1[2][0] = 2093ns;
slave_timing[1][224+6].t_rxd2[0][2] = 2175ns;
slave_timing[1][224+6].t_rxd2[2][0] = 1208ns;
slave_timing[1][224+6].t_rxd2[1][2] = 1834ns;
slave_timing[1][224+6].t_rxd2[2][1] = 1558ns;

slave_timing[1][224+7].info_corner          = 4;
slave_timing[1][224+7].info_temp__j__       = -40;
slave_timing[1][224+7].info_i__quite_rec__  = 0.006000000;
slave_timing[1][224+7].info_dtr__ib__       = 1;
slave_timing[1][224+7].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+7].info_i__max_slave__  = 0.025000000;
slave_timing[1][224+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][224+7].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+7].t_rxd1[0][1] = 1739ns;
slave_timing[1][224+7].t_rxd1[1][0] = 1766ns;
slave_timing[1][224+7].t_rxd1[0][2] = 1312ns;
slave_timing[1][224+7].t_rxd1[2][0] = 2129ns;
slave_timing[1][224+7].t_rxd2[0][2] = 2025ns;
slave_timing[1][224+7].t_rxd2[2][0] = 1302ns;
slave_timing[1][224+7].t_rxd2[1][2] = 1633ns;
slave_timing[1][224+7].t_rxd2[2][1] = 1735ns;

slave_timing[1][224+8].info_corner          = 4;
slave_timing[1][224+8].info_temp__j__       = -40;
slave_timing[1][224+8].info_i__quite_rec__  = 0.003000000;
slave_timing[1][224+8].info_dtr__ib__       = -1;
slave_timing[1][224+8].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+8].info_i__max_slave__  = 0.023000000;
slave_timing[1][224+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][224+8].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+8].t_rxd1[0][1] = 1693ns;
slave_timing[1][224+8].t_rxd1[1][0] = 1691ns;
slave_timing[1][224+8].t_rxd1[0][2] = 1270ns;
slave_timing[1][224+8].t_rxd1[2][0] = 2064ns;
slave_timing[1][224+8].t_rxd2[0][2] = 2049ns;
slave_timing[1][224+8].t_rxd2[2][0] = 1261ns;
slave_timing[1][224+8].t_rxd2[1][2] = 1680ns;
slave_timing[1][224+8].t_rxd2[2][1] = 1672ns;

slave_timing[1][224+9].info_corner          = 4;
slave_timing[1][224+9].info_temp__j__       = -40;
slave_timing[1][224+9].info_i__quite_rec__  = 0.003000000;
slave_timing[1][224+9].info_dtr__ib__       = -1;
slave_timing[1][224+9].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+9].info_i__max_slave__  = 0.025000000;
slave_timing[1][224+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][224+9].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+9].t_rxd1[0][1] = 1627ns;
slave_timing[1][224+9].t_rxd1[1][0] = 1741ns;
slave_timing[1][224+9].t_rxd1[0][2] = 1220ns;
slave_timing[1][224+9].t_rxd1[2][0] = 2101ns;
slave_timing[1][224+9].t_rxd2[0][2] = 1910ns;
slave_timing[1][224+9].t_rxd2[2][0] = 1346ns;
slave_timing[1][224+9].t_rxd2[1][2] = 1500ns;
slave_timing[1][224+9].t_rxd2[2][1] = 1846ns;

slave_timing[1][224+10].info_corner          = 4;
slave_timing[1][224+10].info_temp__j__       = -40;
slave_timing[1][224+10].info_i__quite_rec__  = 0.003000000;
slave_timing[1][224+10].info_dtr__ib__       = 1;
slave_timing[1][224+10].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+10].info_i__max_slave__  = 0.023000000;
slave_timing[1][224+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][224+10].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+10].t_rxd1[0][1] = 1732ns;
slave_timing[1][224+10].t_rxd1[1][0] = 1654ns;
slave_timing[1][224+10].t_rxd1[0][2] = 1276ns;
slave_timing[1][224+10].t_rxd1[2][0] = 2035ns;
slave_timing[1][224+10].t_rxd2[0][2] = 2126ns;
slave_timing[1][224+10].t_rxd2[2][0] = 1197ns;
slave_timing[1][224+10].t_rxd2[1][2] = 1814ns;
slave_timing[1][224+10].t_rxd2[2][1] = 1554ns;

slave_timing[1][224+11].info_corner          = 4;
slave_timing[1][224+11].info_temp__j__       = -40;
slave_timing[1][224+11].info_i__quite_rec__  = 0.003000000;
slave_timing[1][224+11].info_dtr__ib__       = 1;
slave_timing[1][224+11].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+11].info_i__max_slave__  = 0.025000000;
slave_timing[1][224+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][224+11].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+11].t_rxd1[0][1] = 1665ns;
slave_timing[1][224+11].t_rxd1[1][0] = 1706ns;
slave_timing[1][224+11].t_rxd1[0][2] = 1252ns;
slave_timing[1][224+11].t_rxd1[2][0] = 2073ns;
slave_timing[1][224+11].t_rxd2[0][2] = 2000ns;
slave_timing[1][224+11].t_rxd2[2][0] = 1290ns;
slave_timing[1][224+11].t_rxd2[1][2] = 1612ns;
slave_timing[1][224+11].t_rxd2[2][1] = 1729ns;

slave_timing[1][224+12].info_corner          = 4;
slave_timing[1][224+12].info_temp__j__       = -40;
slave_timing[1][224+12].info_i__quite_rec__  = 0.003000000;
slave_timing[1][224+12].info_dtr__ib__       = -1;
slave_timing[1][224+12].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+12].info_i__max_slave__  = 0.023000000;
slave_timing[1][224+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][224+12].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+12].t_rxd1[0][1] = 1771ns;
slave_timing[1][224+12].t_rxd1[1][0] = 1758ns;
slave_timing[1][224+12].t_rxd1[0][2] = 1335ns;
slave_timing[1][224+12].t_rxd1[2][0] = 2133ns;
slave_timing[1][224+12].t_rxd2[0][2] = 2069ns;
slave_timing[1][224+12].t_rxd2[2][0] = 1276ns;
slave_timing[1][224+12].t_rxd2[1][2] = 1715ns;
slave_timing[1][224+12].t_rxd2[2][1] = 1654ns;

slave_timing[1][224+13].info_corner          = 4;
slave_timing[1][224+13].info_temp__j__       = -40;
slave_timing[1][224+13].info_i__quite_rec__  = 0.003000000;
slave_timing[1][224+13].info_dtr__ib__       = -1;
slave_timing[1][224+13].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+13].info_i__max_slave__  = 0.025000000;
slave_timing[1][224+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][224+13].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+13].t_rxd1[0][1] = 1704ns;
slave_timing[1][224+13].t_rxd1[1][0] = 1812ns;
slave_timing[1][224+13].t_rxd1[0][2] = 1296ns;
slave_timing[1][224+13].t_rxd1[2][0] = 2168ns;
slave_timing[1][224+13].t_rxd2[0][2] = 1944ns;
slave_timing[1][224+13].t_rxd2[2][0] = 1360ns;
slave_timing[1][224+13].t_rxd2[1][2] = 1511ns;
slave_timing[1][224+13].t_rxd2[2][1] = 1855ns;

slave_timing[1][224+14].info_corner          = 4;
slave_timing[1][224+14].info_temp__j__       = -40;
slave_timing[1][224+14].info_i__quite_rec__  = 0.003000000;
slave_timing[1][224+14].info_dtr__ib__       = 1;
slave_timing[1][224+14].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+14].info_i__max_slave__  = 0.023000000;
slave_timing[1][224+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][224+14].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+14].t_rxd1[0][1] = 1809ns;
slave_timing[1][224+14].t_rxd1[1][0] = 1721ns;
slave_timing[1][224+14].t_rxd1[0][2] = 1350ns;
slave_timing[1][224+14].t_rxd1[2][0] = 2101ns;
slave_timing[1][224+14].t_rxd2[0][2] = 2167ns;
slave_timing[1][224+14].t_rxd2[2][0] = 1212ns;
slave_timing[1][224+14].t_rxd2[1][2] = 1822ns;
slave_timing[1][224+14].t_rxd2[2][1] = 1564ns;

slave_timing[1][224+15].info_corner          = 4;
slave_timing[1][224+15].info_temp__j__       = -40;
slave_timing[1][224+15].info_i__quite_rec__  = 0.003000000;
slave_timing[1][224+15].info_dtr__ib__       = 1;
slave_timing[1][224+15].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+15].info_i__max_slave__  = 0.025000000;
slave_timing[1][224+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][224+15].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+15].t_rxd1[0][1] = 1735ns;
slave_timing[1][224+15].t_rxd1[1][0] = 1773ns;
slave_timing[1][224+15].t_rxd1[0][2] = 1310ns;
slave_timing[1][224+15].t_rxd1[2][0] = 2137ns;
slave_timing[1][224+15].t_rxd2[0][2] = 2018ns;
slave_timing[1][224+15].t_rxd2[2][0] = 1304ns;
slave_timing[1][224+15].t_rxd2[1][2] = 1624ns;
slave_timing[1][224+15].t_rxd2[2][1] = 1739ns;

slave_timing[1][224+16].info_corner          = 4;
slave_timing[1][224+16].info_temp__j__       = -40;
slave_timing[1][224+16].info_i__quite_rec__  = 0.000000000;
slave_timing[1][224+16].info_dtr__ib__       = -1;
slave_timing[1][224+16].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+16].info_i__max_slave__  = 0.023000000;
slave_timing[1][224+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][224+16].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+16].t_rxd1[0][1] = 1707ns;
slave_timing[1][224+16].t_rxd1[1][0] = 1678ns;
slave_timing[1][224+16].t_rxd1[0][2] = 1262ns;
slave_timing[1][224+16].t_rxd1[2][0] = 2054ns;
slave_timing[1][224+16].t_rxd2[0][2] = 2040ns;
slave_timing[1][224+16].t_rxd2[2][0] = 1258ns;
slave_timing[1][224+16].t_rxd2[1][2] = 1695ns;
slave_timing[1][224+16].t_rxd2[2][1] = 1660ns;

slave_timing[1][224+17].info_corner          = 4;
slave_timing[1][224+17].info_temp__j__       = -40;
slave_timing[1][224+17].info_i__quite_rec__  = 0.000000000;
slave_timing[1][224+17].info_dtr__ib__       = -1;
slave_timing[1][224+17].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+17].info_i__max_slave__  = 0.025000000;
slave_timing[1][224+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][224+17].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+17].t_rxd1[0][1] = 1639ns;
slave_timing[1][224+17].t_rxd1[1][0] = 1730ns;
slave_timing[1][224+17].t_rxd1[0][2] = 1229ns;
slave_timing[1][224+17].t_rxd1[2][0] = 2091ns;
slave_timing[1][224+17].t_rxd2[0][2] = 1918ns;
slave_timing[1][224+17].t_rxd2[2][0] = 1343ns;
slave_timing[1][224+17].t_rxd2[1][2] = 1512ns;
slave_timing[1][224+17].t_rxd2[2][1] = 1838ns;

slave_timing[1][224+18].info_corner          = 4;
slave_timing[1][224+18].info_temp__j__       = -40;
slave_timing[1][224+18].info_i__quite_rec__  = 0.000000000;
slave_timing[1][224+18].info_dtr__ib__       = 1;
slave_timing[1][224+18].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+18].info_i__max_slave__  = 0.023000000;
slave_timing[1][224+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][224+18].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+18].t_rxd1[0][1] = 1725ns;
slave_timing[1][224+18].t_rxd1[1][0] = 1668ns;
slave_timing[1][224+18].t_rxd1[0][2] = 1287ns;
slave_timing[1][224+18].t_rxd1[2][0] = 2044ns;
slave_timing[1][224+18].t_rxd2[0][2] = 2140ns;
slave_timing[1][224+18].t_rxd2[2][0] = 1202ns;
slave_timing[1][224+18].t_rxd2[1][2] = 1819ns;
slave_timing[1][224+18].t_rxd2[2][1] = 1540ns;

slave_timing[1][224+19].info_corner          = 4;
slave_timing[1][224+19].info_temp__j__       = -40;
slave_timing[1][224+19].info_i__quite_rec__  = 0.000000000;
slave_timing[1][224+19].info_dtr__ib__       = 1;
slave_timing[1][224+19].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+19].info_i__max_slave__  = 0.025000000;
slave_timing[1][224+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][224+19].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+19].t_rxd1[0][1] = 1654ns;
slave_timing[1][224+19].t_rxd1[1][0] = 1721ns;
slave_timing[1][224+19].t_rxd1[0][2] = 1249ns;
slave_timing[1][224+19].t_rxd1[2][0] = 2082ns;
slave_timing[1][224+19].t_rxd2[0][2] = 1993ns;
slave_timing[1][224+19].t_rxd2[2][0] = 1295ns;
slave_timing[1][224+19].t_rxd2[1][2] = 1602ns;
slave_timing[1][224+19].t_rxd2[2][1] = 1735ns;

slave_timing[1][224+20].info_corner          = 4;
slave_timing[1][224+20].info_temp__j__       = -40;
slave_timing[1][224+20].info_i__quite_rec__  = 0.000000000;
slave_timing[1][224+20].info_dtr__ib__       = -1;
slave_timing[1][224+20].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+20].info_i__max_slave__  = 0.023000000;
slave_timing[1][224+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][224+20].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+20].t_rxd1[0][1] = 1790ns;
slave_timing[1][224+20].t_rxd1[1][0] = 1749ns;
slave_timing[1][224+20].t_rxd1[0][2] = 1330ns;
slave_timing[1][224+20].t_rxd1[2][0] = 2122ns;
slave_timing[1][224+20].t_rxd2[0][2] = 2060ns;
slave_timing[1][224+20].t_rxd2[2][0] = 1271ns;
slave_timing[1][224+20].t_rxd2[1][2] = 1704ns;
slave_timing[1][224+20].t_rxd2[2][1] = 1671ns;

slave_timing[1][224+21].info_corner          = 4;
slave_timing[1][224+21].info_temp__j__       = -40;
slave_timing[1][224+21].info_i__quite_rec__  = 0.000000000;
slave_timing[1][224+21].info_dtr__ib__       = -1;
slave_timing[1][224+21].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+21].info_i__max_slave__  = 0.025000000;
slave_timing[1][224+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][224+21].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+21].t_rxd1[0][1] = 1720ns;
slave_timing[1][224+21].t_rxd1[1][0] = 1800ns;
slave_timing[1][224+21].t_rxd1[0][2] = 1292ns;
slave_timing[1][224+21].t_rxd1[2][0] = 2159ns;
slave_timing[1][224+21].t_rxd2[0][2] = 1938ns;
slave_timing[1][224+21].t_rxd2[2][0] = 1356ns;
slave_timing[1][224+21].t_rxd2[1][2] = 1521ns;
slave_timing[1][224+21].t_rxd2[2][1] = 1845ns;

slave_timing[1][224+22].info_corner          = 4;
slave_timing[1][224+22].info_temp__j__       = -40;
slave_timing[1][224+22].info_i__quite_rec__  = 0.000000000;
slave_timing[1][224+22].info_dtr__ib__       = 1;
slave_timing[1][224+22].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+22].info_i__max_slave__  = 0.023000000;
slave_timing[1][224+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][224+22].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+22].t_rxd1[0][1] = 1833ns;
slave_timing[1][224+22].t_rxd1[1][0] = 1705ns;
slave_timing[1][224+22].t_rxd1[0][2] = 1346ns;
slave_timing[1][224+22].t_rxd1[2][0] = 2110ns;
slave_timing[1][224+22].t_rxd2[0][2] = 2156ns;
slave_timing[1][224+22].t_rxd2[2][0] = 1216ns;
slave_timing[1][224+22].t_rxd2[1][2] = 1839ns;
slave_timing[1][224+22].t_rxd2[2][1] = 1547ns;

slave_timing[1][224+23].info_corner          = 4;
slave_timing[1][224+23].info_temp__j__       = -40;
slave_timing[1][224+23].info_i__quite_rec__  = 0.000000000;
slave_timing[1][224+23].info_dtr__ib__       = 1;
slave_timing[1][224+23].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+23].info_i__max_slave__  = 0.025000000;
slave_timing[1][224+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][224+23].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+23].t_rxd1[0][1] = 1730ns;
slave_timing[1][224+23].t_rxd1[1][0] = 1785ns;
slave_timing[1][224+23].t_rxd1[0][2] = 1309ns;
slave_timing[1][224+23].t_rxd1[2][0] = 2146ns;
slave_timing[1][224+23].t_rxd2[0][2] = 2010ns;
slave_timing[1][224+23].t_rxd2[2][0] = 1305ns;
slave_timing[1][224+23].t_rxd2[1][2] = 1615ns;
slave_timing[1][224+23].t_rxd2[2][1] = 1746ns;

slave_timing[1][224+24].info_corner          = 4;
slave_timing[1][224+24].info_temp__j__       = -40;
slave_timing[1][224+24].info_i__quite_rec__  = 0.040000000;
slave_timing[1][224+24].info_dtr__ib__       = -1;
slave_timing[1][224+24].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+24].info_i__max_slave__  = 0.023000000;
slave_timing[1][224+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][224+24].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+24].t_rxd1[0][1] = 1675ns;
slave_timing[1][224+24].t_rxd1[1][0] = 1687ns;
slave_timing[1][224+24].t_rxd1[0][2] = 1257ns;
slave_timing[1][224+24].t_rxd1[2][0] = 2056ns;
slave_timing[1][224+24].t_rxd2[0][2] = 2044ns;
slave_timing[1][224+24].t_rxd2[2][0] = 1266ns;
slave_timing[1][224+24].t_rxd2[1][2] = 1701ns;
slave_timing[1][224+24].t_rxd2[2][1] = 1654ns;

slave_timing[1][224+25].info_corner          = 4;
slave_timing[1][224+25].info_temp__j__       = -40;
slave_timing[1][224+25].info_i__quite_rec__  = 0.040000000;
slave_timing[1][224+25].info_dtr__ib__       = -1;
slave_timing[1][224+25].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+25].info_i__max_slave__  = 0.025000000;
slave_timing[1][224+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][224+25].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+25].t_rxd1[0][1] = 1611ns;
slave_timing[1][224+25].t_rxd1[1][0] = 1739ns;
slave_timing[1][224+25].t_rxd1[0][2] = 1224ns;
slave_timing[1][224+25].t_rxd1[2][0] = 2092ns;
slave_timing[1][224+25].t_rxd2[0][2] = 1920ns;
slave_timing[1][224+25].t_rxd2[2][0] = 1349ns;
slave_timing[1][224+25].t_rxd2[1][2] = 1495ns;
slave_timing[1][224+25].t_rxd2[2][1] = 1856ns;

slave_timing[1][224+26].info_corner          = 4;
slave_timing[1][224+26].info_temp__j__       = -40;
slave_timing[1][224+26].info_i__quite_rec__  = 0.040000000;
slave_timing[1][224+26].info_dtr__ib__       = 1;
slave_timing[1][224+26].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+26].info_i__max_slave__  = 0.023000000;
slave_timing[1][224+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][224+26].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+26].t_rxd1[0][1] = 1728ns;
slave_timing[1][224+26].t_rxd1[1][0] = 1645ns;
slave_timing[1][224+26].t_rxd1[0][2] = 1286ns;
slave_timing[1][224+26].t_rxd1[2][0] = 2026ns;
slave_timing[1][224+26].t_rxd2[0][2] = 2150ns;
slave_timing[1][224+26].t_rxd2[2][0] = 1198ns;
slave_timing[1][224+26].t_rxd2[1][2] = 1820ns;
slave_timing[1][224+26].t_rxd2[2][1] = 1554ns;

slave_timing[1][224+27].info_corner          = 4;
slave_timing[1][224+27].info_temp__j__       = -40;
slave_timing[1][224+27].info_i__quite_rec__  = 0.040000000;
slave_timing[1][224+27].info_dtr__ib__       = 1;
slave_timing[1][224+27].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+27].info_i__max_slave__  = 0.025000000;
slave_timing[1][224+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][224+27].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+27].t_rxd1[0][1] = 1658ns;
slave_timing[1][224+27].t_rxd1[1][0] = 1698ns;
slave_timing[1][224+27].t_rxd1[0][2] = 1248ns;
slave_timing[1][224+27].t_rxd1[2][0] = 2063ns;
slave_timing[1][224+27].t_rxd2[0][2] = 2002ns;
slave_timing[1][224+27].t_rxd2[2][0] = 1289ns;
slave_timing[1][224+27].t_rxd2[1][2] = 1619ns;
slave_timing[1][224+27].t_rxd2[2][1] = 1728ns;

slave_timing[1][224+28].info_corner          = 4;
slave_timing[1][224+28].info_temp__j__       = -40;
slave_timing[1][224+28].info_i__quite_rec__  = 0.040000000;
slave_timing[1][224+28].info_dtr__ib__       = -1;
slave_timing[1][224+28].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+28].info_i__max_slave__  = 0.023000000;
slave_timing[1][224+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][224+28].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+28].t_rxd1[0][1] = 1714ns;
slave_timing[1][224+28].t_rxd1[1][0] = 1721ns;
slave_timing[1][224+28].t_rxd1[0][2] = 1293ns;
slave_timing[1][224+28].t_rxd1[2][0] = 2088ns;
slave_timing[1][224+28].t_rxd2[0][2] = 2061ns;
slave_timing[1][224+28].t_rxd2[2][0] = 1281ns;
slave_timing[1][224+28].t_rxd2[1][2] = 1694ns;
slave_timing[1][224+28].t_rxd2[2][1] = 1671ns;

slave_timing[1][224+29].info_corner          = 4;
slave_timing[1][224+29].info_temp__j__       = -40;
slave_timing[1][224+29].info_i__quite_rec__  = 0.040000000;
slave_timing[1][224+29].info_dtr__ib__       = -1;
slave_timing[1][224+29].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+29].info_i__max_slave__  = 0.025000000;
slave_timing[1][224+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][224+29].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+29].t_rxd1[0][1] = 1647ns;
slave_timing[1][224+29].t_rxd1[1][0] = 1775ns;
slave_timing[1][224+29].t_rxd1[0][2] = 1258ns;
slave_timing[1][224+29].t_rxd1[2][0] = 2124ns;
slave_timing[1][224+29].t_rxd2[0][2] = 1941ns;
slave_timing[1][224+29].t_rxd2[2][0] = 1366ns;
slave_timing[1][224+29].t_rxd2[1][2] = 1518ns;
slave_timing[1][224+29].t_rxd2[2][1] = 1863ns;

slave_timing[1][224+30].info_corner          = 4;
slave_timing[1][224+30].info_temp__j__       = -40;
slave_timing[1][224+30].info_i__quite_rec__  = 0.040000000;
slave_timing[1][224+30].info_dtr__ib__       = 1;
slave_timing[1][224+30].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+30].info_i__max_slave__  = 0.023000000;
slave_timing[1][224+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][224+30].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+30].t_rxd1[0][1] = 1764ns;
slave_timing[1][224+30].t_rxd1[1][0] = 1679ns;
slave_timing[1][224+30].t_rxd1[0][2] = 1320ns;
slave_timing[1][224+30].t_rxd1[2][0] = 2056ns;
slave_timing[1][224+30].t_rxd2[0][2] = 2164ns;
slave_timing[1][224+30].t_rxd2[2][0] = 1214ns;
slave_timing[1][224+30].t_rxd2[1][2] = 1836ns;
slave_timing[1][224+30].t_rxd2[2][1] = 1565ns;

slave_timing[1][224+31].info_corner          = 4;
slave_timing[1][224+31].info_temp__j__       = -40;
slave_timing[1][224+31].info_i__quite_rec__  = 0.040000000;
slave_timing[1][224+31].info_dtr__ib__       = 1;
slave_timing[1][224+31].info_i__offset_rec__ = 0.000000000;
slave_timing[1][224+31].info_i__max_slave__  = 0.025000000;
slave_timing[1][224+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][224+31].info_r__dsi_bus__    = 5.000;

slave_timing[1][224+31].t_rxd1[0][1] = 1693ns;
slave_timing[1][224+31].t_rxd1[1][0] = 1732ns;
slave_timing[1][224+31].t_rxd1[0][2] = 1281ns;
slave_timing[1][224+31].t_rxd1[2][0] = 2092ns;
slave_timing[1][224+31].t_rxd2[0][2] = 2018ns;
slave_timing[1][224+31].t_rxd2[2][0] = 1306ns;
slave_timing[1][224+31].t_rxd2[1][2] = 1638ns;
slave_timing[1][224+31].t_rxd2[2][1] = 1738ns;

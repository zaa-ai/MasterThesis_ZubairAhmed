
slave_timing[3][128+0].info_corner          = 1;
slave_timing[3][128+0].info_temp__j__       = -40;
slave_timing[3][128+0].info_i__quite_rec__  = 0.006000000;
slave_timing[3][128+0].info_dtr__ib__       = -1;
slave_timing[3][128+0].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+0].info_i__max_slave__  = 0.023000000;
slave_timing[3][128+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][128+0].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+0].t_rxd1[0][1] = 2681ns;
slave_timing[3][128+0].t_rxd1[1][0] = 2717ns;
slave_timing[3][128+0].t_rxd1[0][2] = 1983ns;
slave_timing[3][128+0].t_rxd1[2][0] = 3311ns;
slave_timing[3][128+0].t_rxd2[0][2] = 3248ns;
slave_timing[3][128+0].t_rxd2[2][0] = 2029ns;
slave_timing[3][128+0].t_rxd2[1][2] = 2656ns;
slave_timing[3][128+0].t_rxd2[2][1] = 2710ns;

slave_timing[3][128+1].info_corner          = 1;
slave_timing[3][128+1].info_temp__j__       = -40;
slave_timing[3][128+1].info_i__quite_rec__  = 0.006000000;
slave_timing[3][128+1].info_dtr__ib__       = -1;
slave_timing[3][128+1].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+1].info_i__max_slave__  = 0.025000000;
slave_timing[3][128+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][128+1].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+1].t_rxd1[0][1] = 2579ns;
slave_timing[3][128+1].t_rxd1[1][0] = 2799ns;
slave_timing[3][128+1].t_rxd1[0][2] = 1947ns;
slave_timing[3][128+1].t_rxd1[2][0] = 3362ns;
slave_timing[3][128+1].t_rxd2[0][2] = 3071ns;
slave_timing[3][128+1].t_rxd2[2][0] = 2174ns;
slave_timing[3][128+1].t_rxd2[1][2] = 2379ns;
slave_timing[3][128+1].t_rxd2[2][1] = 2999ns;

slave_timing[3][128+2].info_corner          = 1;
slave_timing[3][128+2].info_temp__j__       = -40;
slave_timing[3][128+2].info_i__quite_rec__  = 0.006000000;
slave_timing[3][128+2].info_dtr__ib__       = 1;
slave_timing[3][128+2].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+2].info_i__max_slave__  = 0.023000000;
slave_timing[3][128+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][128+2].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+2].t_rxd1[0][1] = 2792ns;
slave_timing[3][128+2].t_rxd1[1][0] = 2639ns;
slave_timing[3][128+2].t_rxd1[0][2] = 2069ns;
slave_timing[3][128+2].t_rxd1[2][0] = 3256ns;
slave_timing[3][128+2].t_rxd2[0][2] = 3455ns;
slave_timing[3][128+2].t_rxd2[2][0] = 1874ns;
slave_timing[3][128+2].t_rxd2[1][2] = 2951ns;
slave_timing[3][128+2].t_rxd2[2][1] = 2463ns;

slave_timing[3][128+3].info_corner          = 1;
slave_timing[3][128+3].info_temp__j__       = -40;
slave_timing[3][128+3].info_i__quite_rec__  = 0.006000000;
slave_timing[3][128+3].info_dtr__ib__       = 1;
slave_timing[3][128+3].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+3].info_i__max_slave__  = 0.025000000;
slave_timing[3][128+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][128+3].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+3].t_rxd1[0][1] = 2676ns;
slave_timing[3][128+3].t_rxd1[1][0] = 2722ns;
slave_timing[3][128+3].t_rxd1[0][2] = 2003ns;
slave_timing[3][128+3].t_rxd1[2][0] = 3311ns;
slave_timing[3][128+3].t_rxd2[0][2] = 3229ns;
slave_timing[3][128+3].t_rxd2[2][0] = 2045ns;
slave_timing[3][128+3].t_rxd2[1][2] = 2661ns;
slave_timing[3][128+3].t_rxd2[2][1] = 2708ns;

slave_timing[3][128+4].info_corner          = 1;
slave_timing[3][128+4].info_temp__j__       = -40;
slave_timing[3][128+4].info_i__quite_rec__  = 0.006000000;
slave_timing[3][128+4].info_dtr__ib__       = -1;
slave_timing[3][128+4].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+4].info_i__max_slave__  = 0.023000000;
slave_timing[3][128+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][128+4].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+4].t_rxd1[0][1] = 2756ns;
slave_timing[3][128+4].t_rxd1[1][0] = 2789ns;
slave_timing[3][128+4].t_rxd1[0][2] = 2076ns;
slave_timing[3][128+4].t_rxd1[2][0] = 3380ns;
slave_timing[3][128+4].t_rxd2[0][2] = 3268ns;
slave_timing[3][128+4].t_rxd2[2][0] = 2043ns;
slave_timing[3][128+4].t_rxd2[1][2] = 2671ns;
slave_timing[3][128+4].t_rxd2[2][1] = 2727ns;

slave_timing[3][128+5].info_corner          = 1;
slave_timing[3][128+5].info_temp__j__       = -40;
slave_timing[3][128+5].info_i__quite_rec__  = 0.006000000;
slave_timing[3][128+5].info_dtr__ib__       = -1;
slave_timing[3][128+5].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+5].info_i__max_slave__  = 0.025000000;
slave_timing[3][128+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][128+5].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+5].t_rxd1[0][1] = 2655ns;
slave_timing[3][128+5].t_rxd1[1][0] = 2873ns;
slave_timing[3][128+5].t_rxd1[0][2] = 2017ns;
slave_timing[3][128+5].t_rxd1[2][0] = 3433ns;
slave_timing[3][128+5].t_rxd2[0][2] = 3086ns;
slave_timing[3][128+5].t_rxd2[2][0] = 2189ns;
slave_timing[3][128+5].t_rxd2[1][2] = 2381ns;
slave_timing[3][128+5].t_rxd2[2][1] = 3009ns;

slave_timing[3][128+6].info_corner          = 1;
slave_timing[3][128+6].info_temp__j__       = -40;
slave_timing[3][128+6].info_i__quite_rec__  = 0.006000000;
slave_timing[3][128+6].info_dtr__ib__       = 1;
slave_timing[3][128+6].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+6].info_i__max_slave__  = 0.023000000;
slave_timing[3][128+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][128+6].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+6].t_rxd1[0][1] = 2860ns;
slave_timing[3][128+6].t_rxd1[1][0] = 2703ns;
slave_timing[3][128+6].t_rxd1[0][2] = 2134ns;
slave_timing[3][128+6].t_rxd1[2][0] = 3327ns;
slave_timing[3][128+6].t_rxd2[0][2] = 3469ns;
slave_timing[3][128+6].t_rxd2[2][0] = 1889ns;
slave_timing[3][128+6].t_rxd2[1][2] = 2959ns;
slave_timing[3][128+6].t_rxd2[2][1] = 2439ns;

slave_timing[3][128+7].info_corner          = 1;
slave_timing[3][128+7].info_temp__j__       = -40;
slave_timing[3][128+7].info_i__quite_rec__  = 0.006000000;
slave_timing[3][128+7].info_dtr__ib__       = 1;
slave_timing[3][128+7].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+7].info_i__max_slave__  = 0.025000000;
slave_timing[3][128+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][128+7].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+7].t_rxd1[0][1] = 2750ns;
slave_timing[3][128+7].t_rxd1[1][0] = 2795ns;
slave_timing[3][128+7].t_rxd1[0][2] = 2067ns;
slave_timing[3][128+7].t_rxd1[2][0] = 3380ns;
slave_timing[3][128+7].t_rxd2[0][2] = 3243ns;
slave_timing[3][128+7].t_rxd2[2][0] = 2060ns;
slave_timing[3][128+7].t_rxd2[1][2] = 2633ns;
slave_timing[3][128+7].t_rxd2[2][1] = 2715ns;

slave_timing[3][128+8].info_corner          = 1;
slave_timing[3][128+8].info_temp__j__       = -40;
slave_timing[3][128+8].info_i__quite_rec__  = 0.003000000;
slave_timing[3][128+8].info_dtr__ib__       = -1;
slave_timing[3][128+8].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+8].info_i__max_slave__  = 0.023000000;
slave_timing[3][128+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][128+8].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+8].t_rxd1[0][1] = 2710ns;
slave_timing[3][128+8].t_rxd1[1][0] = 2688ns;
slave_timing[3][128+8].t_rxd1[0][2] = 2025ns;
slave_timing[3][128+8].t_rxd1[2][0] = 3293ns;
slave_timing[3][128+8].t_rxd2[0][2] = 3272ns;
slave_timing[3][128+8].t_rxd2[2][0] = 2015ns;
slave_timing[3][128+8].t_rxd2[1][2] = 2683ns;
slave_timing[3][128+8].t_rxd2[2][1] = 2654ns;

slave_timing[3][128+9].info_corner          = 1;
slave_timing[3][128+9].info_temp__j__       = -40;
slave_timing[3][128+9].info_i__quite_rec__  = 0.003000000;
slave_timing[3][128+9].info_dtr__ib__       = -1;
slave_timing[3][128+9].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+9].info_i__max_slave__  = 0.025000000;
slave_timing[3][128+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][128+9].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+9].t_rxd1[0][1] = 2612ns;
slave_timing[3][128+9].t_rxd1[1][0] = 2775ns;
slave_timing[3][128+9].t_rxd1[0][2] = 1961ns;
slave_timing[3][128+9].t_rxd1[2][0] = 3346ns;
slave_timing[3][128+9].t_rxd2[0][2] = 3083ns;
slave_timing[3][128+9].t_rxd2[2][0] = 2164ns;
slave_timing[3][128+9].t_rxd2[1][2] = 2402ns;
slave_timing[3][128+9].t_rxd2[2][1] = 2976ns;

slave_timing[3][128+10].info_corner          = 1;
slave_timing[3][128+10].info_temp__j__       = -40;
slave_timing[3][128+10].info_i__quite_rec__  = 0.003000000;
slave_timing[3][128+10].info_dtr__ib__       = 1;
slave_timing[3][128+10].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+10].info_i__max_slave__  = 0.023000000;
slave_timing[3][128+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][128+10].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+10].t_rxd1[0][1] = 2819ns;
slave_timing[3][128+10].t_rxd1[1][0] = 2608ns;
slave_timing[3][128+10].t_rxd1[0][2] = 2081ns;
slave_timing[3][128+10].t_rxd1[2][0] = 3236ns;
slave_timing[3][128+10].t_rxd2[0][2] = 3480ns;
slave_timing[3][128+10].t_rxd2[2][0] = 1861ns;
slave_timing[3][128+10].t_rxd2[1][2] = 2970ns;
slave_timing[3][128+10].t_rxd2[2][1] = 2446ns;

slave_timing[3][128+11].info_corner          = 1;
slave_timing[3][128+11].info_temp__j__       = -40;
slave_timing[3][128+11].info_i__quite_rec__  = 0.003000000;
slave_timing[3][128+11].info_dtr__ib__       = 1;
slave_timing[3][128+11].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+11].info_i__max_slave__  = 0.025000000;
slave_timing[3][128+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][128+11].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+11].t_rxd1[0][1] = 2703ns;
slave_timing[3][128+11].t_rxd1[1][0] = 2694ns;
slave_timing[3][128+11].t_rxd1[0][2] = 2014ns;
slave_timing[3][128+11].t_rxd1[2][0] = 3291ns;
slave_timing[3][128+11].t_rxd2[0][2] = 3251ns;
slave_timing[3][128+11].t_rxd2[2][0] = 2031ns;
slave_timing[3][128+11].t_rxd2[1][2] = 2644ns;
slave_timing[3][128+11].t_rxd2[2][1] = 2730ns;

slave_timing[3][128+12].info_corner          = 1;
slave_timing[3][128+12].info_temp__j__       = -40;
slave_timing[3][128+12].info_i__quite_rec__  = 0.003000000;
slave_timing[3][128+12].info_dtr__ib__       = -1;
slave_timing[3][128+12].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+12].info_i__max_slave__  = 0.023000000;
slave_timing[3][128+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][128+12].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+12].t_rxd1[0][1] = 2784ns;
slave_timing[3][128+12].t_rxd1[1][0] = 2764ns;
slave_timing[3][128+12].t_rxd1[0][2] = 2090ns;
slave_timing[3][128+12].t_rxd1[2][0] = 3362ns;
slave_timing[3][128+12].t_rxd2[0][2] = 3282ns;
slave_timing[3][128+12].t_rxd2[2][0] = 2033ns;
slave_timing[3][128+12].t_rxd2[1][2] = 2697ns;
slave_timing[3][128+12].t_rxd2[2][1] = 2705ns;

slave_timing[3][128+13].info_corner          = 1;
slave_timing[3][128+13].info_temp__j__       = -40;
slave_timing[3][128+13].info_i__quite_rec__  = 0.003000000;
slave_timing[3][128+13].info_dtr__ib__       = -1;
slave_timing[3][128+13].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+13].info_i__max_slave__  = 0.025000000;
slave_timing[3][128+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][128+13].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+13].t_rxd1[0][1] = 2679ns;
slave_timing[3][128+13].t_rxd1[1][0] = 2847ns;
slave_timing[3][128+13].t_rxd1[0][2] = 2026ns;
slave_timing[3][128+13].t_rxd1[2][0] = 3418ns;
slave_timing[3][128+13].t_rxd2[0][2] = 3093ns;
slave_timing[3][128+13].t_rxd2[2][0] = 2179ns;
slave_timing[3][128+13].t_rxd2[1][2] = 2407ns;
slave_timing[3][128+13].t_rxd2[2][1] = 2988ns;

slave_timing[3][128+14].info_corner          = 1;
slave_timing[3][128+14].info_temp__j__       = -40;
slave_timing[3][128+14].info_i__quite_rec__  = 0.003000000;
slave_timing[3][128+14].info_dtr__ib__       = 1;
slave_timing[3][128+14].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+14].info_i__max_slave__  = 0.023000000;
slave_timing[3][128+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][128+14].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+14].t_rxd1[0][1] = 2893ns;
slave_timing[3][128+14].t_rxd1[1][0] = 2677ns;
slave_timing[3][128+14].t_rxd1[0][2] = 2154ns;
slave_timing[3][128+14].t_rxd1[2][0] = 3305ns;
slave_timing[3][128+14].t_rxd2[0][2] = 3485ns;
slave_timing[3][128+14].t_rxd2[2][0] = 1877ns;
slave_timing[3][128+14].t_rxd2[1][2] = 2983ns;
slave_timing[3][128+14].t_rxd2[2][1] = 2455ns;

slave_timing[3][128+15].info_corner          = 1;
slave_timing[3][128+15].info_temp__j__       = -40;
slave_timing[3][128+15].info_i__quite_rec__  = 0.003000000;
slave_timing[3][128+15].info_dtr__ib__       = 1;
slave_timing[3][128+15].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+15].info_i__max_slave__  = 0.025000000;
slave_timing[3][128+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][128+15].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+15].t_rxd1[0][1] = 2779ns;
slave_timing[3][128+15].t_rxd1[1][0] = 2767ns;
slave_timing[3][128+15].t_rxd1[0][2] = 2086ns;
slave_timing[3][128+15].t_rxd1[2][0] = 3361ns;
slave_timing[3][128+15].t_rxd2[0][2] = 3259ns;
slave_timing[3][128+15].t_rxd2[2][0] = 2052ns;
slave_timing[3][128+15].t_rxd2[1][2] = 2655ns;
slave_timing[3][128+15].t_rxd2[2][1] = 2742ns;

slave_timing[3][128+16].info_corner          = 1;
slave_timing[3][128+16].info_temp__j__       = -40;
slave_timing[3][128+16].info_i__quite_rec__  = 0.000000000;
slave_timing[3][128+16].info_dtr__ib__       = -1;
slave_timing[3][128+16].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+16].info_i__max_slave__  = 0.023000000;
slave_timing[3][128+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][128+16].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+16].t_rxd1[0][1] = 2700ns;
slave_timing[3][128+16].t_rxd1[1][0] = 2706ns;
slave_timing[3][128+16].t_rxd1[0][2] = 2015ns;
slave_timing[3][128+16].t_rxd1[2][0] = 3301ns;
slave_timing[3][128+16].t_rxd2[0][2] = 3261ns;
slave_timing[3][128+16].t_rxd2[2][0] = 2026ns;
slave_timing[3][128+16].t_rxd2[1][2] = 2665ns;
slave_timing[3][128+16].t_rxd2[2][1] = 2712ns;

slave_timing[3][128+17].info_corner          = 1;
slave_timing[3][128+17].info_temp__j__       = -40;
slave_timing[3][128+17].info_i__quite_rec__  = 0.000000000;
slave_timing[3][128+17].info_dtr__ib__       = -1;
slave_timing[3][128+17].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+17].info_i__max_slave__  = 0.025000000;
slave_timing[3][128+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][128+17].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+17].t_rxd1[0][1] = 2595ns;
slave_timing[3][128+17].t_rxd1[1][0] = 2788ns;
slave_timing[3][128+17].t_rxd1[0][2] = 1929ns;
slave_timing[3][128+17].t_rxd1[2][0] = 3354ns;
slave_timing[3][128+17].t_rxd2[0][2] = 3053ns;
slave_timing[3][128+17].t_rxd2[2][0] = 2173ns;
slave_timing[3][128+17].t_rxd2[1][2] = 2382ns;
slave_timing[3][128+17].t_rxd2[2][1] = 2998ns;

slave_timing[3][128+18].info_corner          = 1;
slave_timing[3][128+18].info_temp__j__       = -40;
slave_timing[3][128+18].info_i__quite_rec__  = 0.000000000;
slave_timing[3][128+18].info_dtr__ib__       = 1;
slave_timing[3][128+18].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+18].info_i__max_slave__  = 0.023000000;
slave_timing[3][128+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][128+18].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+18].t_rxd1[0][1] = 2797ns;
slave_timing[3][128+18].t_rxd1[1][0] = 2627ns;
slave_timing[3][128+18].t_rxd1[0][2] = 2072ns;
slave_timing[3][128+18].t_rxd1[2][0] = 3251ns;
slave_timing[3][128+18].t_rxd2[0][2] = 3460ns;
slave_timing[3][128+18].t_rxd2[2][0] = 1871ns;
slave_timing[3][128+18].t_rxd2[1][2] = 2953ns;
slave_timing[3][128+18].t_rxd2[2][1] = 2455ns;

slave_timing[3][128+19].info_corner          = 1;
slave_timing[3][128+19].info_temp__j__       = -40;
slave_timing[3][128+19].info_i__quite_rec__  = 0.000000000;
slave_timing[3][128+19].info_dtr__ib__       = 1;
slave_timing[3][128+19].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+19].info_i__max_slave__  = 0.025000000;
slave_timing[3][128+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][128+19].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+19].t_rxd1[0][1] = 2682ns;
slave_timing[3][128+19].t_rxd1[1][0] = 2712ns;
slave_timing[3][128+19].t_rxd1[0][2] = 2001ns;
slave_timing[3][128+19].t_rxd1[2][0] = 3306ns;
slave_timing[3][128+19].t_rxd2[0][2] = 3232ns;
slave_timing[3][128+19].t_rxd2[2][0] = 2043ns;
slave_timing[3][128+19].t_rxd2[1][2] = 2628ns;
slave_timing[3][128+19].t_rxd2[2][1] = 2741ns;

slave_timing[3][128+20].info_corner          = 1;
slave_timing[3][128+20].info_temp__j__       = -40;
slave_timing[3][128+20].info_i__quite_rec__  = 0.000000000;
slave_timing[3][128+20].info_dtr__ib__       = -1;
slave_timing[3][128+20].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+20].info_i__max_slave__  = 0.023000000;
slave_timing[3][128+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][128+20].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+20].t_rxd1[0][1] = 2769ns;
slave_timing[3][128+20].t_rxd1[1][0] = 2772ns;
slave_timing[3][128+20].t_rxd1[0][2] = 2082ns;
slave_timing[3][128+20].t_rxd1[2][0] = 3368ns;
slave_timing[3][128+20].t_rxd2[0][2] = 3271ns;
slave_timing[3][128+20].t_rxd2[2][0] = 2046ns;
slave_timing[3][128+20].t_rxd2[1][2] = 2679ns;
slave_timing[3][128+20].t_rxd2[2][1] = 2672ns;

slave_timing[3][128+21].info_corner          = 1;
slave_timing[3][128+21].info_temp__j__       = -40;
slave_timing[3][128+21].info_i__quite_rec__  = 0.000000000;
slave_timing[3][128+21].info_dtr__ib__       = -1;
slave_timing[3][128+21].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+21].info_i__max_slave__  = 0.025000000;
slave_timing[3][128+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][128+21].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+21].t_rxd1[0][1] = 2663ns;
slave_timing[3][128+21].t_rxd1[1][0] = 2857ns;
slave_timing[3][128+21].t_rxd1[0][2] = 2018ns;
slave_timing[3][128+21].t_rxd1[2][0] = 3422ns;
slave_timing[3][128+21].t_rxd2[0][2] = 3086ns;
slave_timing[3][128+21].t_rxd2[2][0] = 2188ns;
slave_timing[3][128+21].t_rxd2[1][2] = 2425ns;
slave_timing[3][128+21].t_rxd2[2][1] = 2967ns;

slave_timing[3][128+22].info_corner          = 1;
slave_timing[3][128+22].info_temp__j__       = -40;
slave_timing[3][128+22].info_i__quite_rec__  = 0.000000000;
slave_timing[3][128+22].info_dtr__ib__       = 1;
slave_timing[3][128+22].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+22].info_i__max_slave__  = 0.023000000;
slave_timing[3][128+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][128+22].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+22].t_rxd1[0][1] = 2864ns;
slave_timing[3][128+22].t_rxd1[1][0] = 2695ns;
slave_timing[3][128+22].t_rxd1[0][2] = 2136ns;
slave_timing[3][128+22].t_rxd1[2][0] = 3318ns;
slave_timing[3][128+22].t_rxd2[0][2] = 3468ns;
slave_timing[3][128+22].t_rxd2[2][0] = 1881ns;
slave_timing[3][128+22].t_rxd2[1][2] = 3011ns;
slave_timing[3][128+22].t_rxd2[2][1] = 2426ns;

slave_timing[3][128+23].info_corner          = 1;
slave_timing[3][128+23].info_temp__j__       = -40;
slave_timing[3][128+23].info_i__quite_rec__  = 0.000000000;
slave_timing[3][128+23].info_dtr__ib__       = 1;
slave_timing[3][128+23].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+23].info_i__max_slave__  = 0.025000000;
slave_timing[3][128+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][128+23].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+23].t_rxd1[0][1] = 2752ns;
slave_timing[3][128+23].t_rxd1[1][0] = 2783ns;
slave_timing[3][128+23].t_rxd1[0][2] = 2069ns;
slave_timing[3][128+23].t_rxd1[2][0] = 3375ns;
slave_timing[3][128+23].t_rxd2[0][2] = 3243ns;
slave_timing[3][128+23].t_rxd2[2][0] = 2052ns;
slave_timing[3][128+23].t_rxd2[1][2] = 2637ns;
slave_timing[3][128+23].t_rxd2[2][1] = 2712ns;

slave_timing[3][128+24].info_corner          = 1;
slave_timing[3][128+24].info_temp__j__       = -40;
slave_timing[3][128+24].info_i__quite_rec__  = 0.040000000;
slave_timing[3][128+24].info_dtr__ib__       = -1;
slave_timing[3][128+24].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+24].info_i__max_slave__  = 0.023000000;
slave_timing[3][128+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][128+24].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+24].t_rxd1[0][1] = 2709ns;
slave_timing[3][128+24].t_rxd1[1][0] = 2674ns;
slave_timing[3][128+24].t_rxd1[0][2] = 2021ns;
slave_timing[3][128+24].t_rxd1[2][0] = 3277ns;
slave_timing[3][128+24].t_rxd2[0][2] = 3283ns;
slave_timing[3][128+24].t_rxd2[2][0] = 2018ns;
slave_timing[3][128+24].t_rxd2[1][2] = 2686ns;
slave_timing[3][128+24].t_rxd2[2][1] = 2688ns;

slave_timing[3][128+25].info_corner          = 1;
slave_timing[3][128+25].info_temp__j__       = -40;
slave_timing[3][128+25].info_i__quite_rec__  = 0.040000000;
slave_timing[3][128+25].info_dtr__ib__       = -1;
slave_timing[3][128+25].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+25].info_i__max_slave__  = 0.025000000;
slave_timing[3][128+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][128+25].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+25].t_rxd1[0][1] = 2607ns;
slave_timing[3][128+25].t_rxd1[1][0] = 2758ns;
slave_timing[3][128+25].t_rxd1[0][2] = 1955ns;
slave_timing[3][128+25].t_rxd1[2][0] = 3333ns;
slave_timing[3][128+25].t_rxd2[0][2] = 3087ns;
slave_timing[3][128+25].t_rxd2[2][0] = 2161ns;
slave_timing[3][128+25].t_rxd2[1][2] = 2402ns;
slave_timing[3][128+25].t_rxd2[2][1] = 2974ns;

slave_timing[3][128+26].info_corner          = 1;
slave_timing[3][128+26].info_temp__j__       = -40;
slave_timing[3][128+26].info_i__quite_rec__  = 0.040000000;
slave_timing[3][128+26].info_dtr__ib__       = 1;
slave_timing[3][128+26].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+26].info_i__max_slave__  = 0.023000000;
slave_timing[3][128+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][128+26].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+26].t_rxd1[0][1] = 2782ns;
slave_timing[3][128+26].t_rxd1[1][0] = 2625ns;
slave_timing[3][128+26].t_rxd1[0][2] = 2059ns;
slave_timing[3][128+26].t_rxd1[2][0] = 3246ns;
slave_timing[3][128+26].t_rxd2[0][2] = 3447ns;
slave_timing[3][128+26].t_rxd2[2][0] = 1878ns;
slave_timing[3][128+26].t_rxd2[1][2] = 2942ns;
slave_timing[3][128+26].t_rxd2[2][1] = 2470ns;

slave_timing[3][128+27].info_corner          = 1;
slave_timing[3][128+27].info_temp__j__       = -40;
slave_timing[3][128+27].info_i__quite_rec__  = 0.040000000;
slave_timing[3][128+27].info_dtr__ib__       = 1;
slave_timing[3][128+27].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+27].info_i__max_slave__  = 0.025000000;
slave_timing[3][128+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][128+27].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+27].t_rxd1[0][1] = 2668ns;
slave_timing[3][128+27].t_rxd1[1][0] = 2715ns;
slave_timing[3][128+27].t_rxd1[0][2] = 1995ns;
slave_timing[3][128+27].t_rxd1[2][0] = 3298ns;
slave_timing[3][128+27].t_rxd2[0][2] = 3226ns;
slave_timing[3][128+27].t_rxd2[2][0] = 2045ns;
slave_timing[3][128+27].t_rxd2[1][2] = 2616ns;
slave_timing[3][128+27].t_rxd2[2][1] = 2716ns;

slave_timing[3][128+28].info_corner          = 1;
slave_timing[3][128+28].info_temp__j__       = -40;
slave_timing[3][128+28].info_i__quite_rec__  = 0.040000000;
slave_timing[3][128+28].info_dtr__ib__       = -1;
slave_timing[3][128+28].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+28].info_i__max_slave__  = 0.023000000;
slave_timing[3][128+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][128+28].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+28].t_rxd1[0][1] = 2750ns;
slave_timing[3][128+28].t_rxd1[1][0] = 2713ns;
slave_timing[3][128+28].t_rxd1[0][2] = 2062ns;
slave_timing[3][128+28].t_rxd1[2][0] = 3320ns;
slave_timing[3][128+28].t_rxd2[0][2] = 3288ns;
slave_timing[3][128+28].t_rxd2[2][0] = 2027ns;
slave_timing[3][128+28].t_rxd2[1][2] = 2739ns;
slave_timing[3][128+28].t_rxd2[2][1] = 2658ns;

slave_timing[3][128+29].info_corner          = 1;
slave_timing[3][128+29].info_temp__j__       = -40;
slave_timing[3][128+29].info_i__quite_rec__  = 0.040000000;
slave_timing[3][128+29].info_dtr__ib__       = -1;
slave_timing[3][128+29].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+29].info_i__max_slave__  = 0.025000000;
slave_timing[3][128+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][128+29].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+29].t_rxd1[0][1] = 2650ns;
slave_timing[3][128+29].t_rxd1[1][0] = 2804ns;
slave_timing[3][128+29].t_rxd1[0][2] = 1970ns;
slave_timing[3][128+29].t_rxd1[2][0] = 3376ns;
slave_timing[3][128+29].t_rxd2[0][2] = 3097ns;
slave_timing[3][128+29].t_rxd2[2][0] = 2177ns;
slave_timing[3][128+29].t_rxd2[1][2] = 2415ns;
slave_timing[3][128+29].t_rxd2[2][1] = 2982ns;

slave_timing[3][128+30].info_corner          = 1;
slave_timing[3][128+30].info_temp__j__       = -40;
slave_timing[3][128+30].info_i__quite_rec__  = 0.040000000;
slave_timing[3][128+30].info_dtr__ib__       = 1;
slave_timing[3][128+30].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+30].info_i__max_slave__  = 0.023000000;
slave_timing[3][128+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][128+30].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+30].t_rxd1[0][1] = 2824ns;
slave_timing[3][128+30].t_rxd1[1][0] = 2672ns;
slave_timing[3][128+30].t_rxd1[0][2] = 2098ns;
slave_timing[3][128+30].t_rxd1[2][0] = 3291ns;
slave_timing[3][128+30].t_rxd2[0][2] = 3461ns;
slave_timing[3][128+30].t_rxd2[2][0] = 1888ns;
slave_timing[3][128+30].t_rxd2[1][2] = 2946ns;
slave_timing[3][128+30].t_rxd2[2][1] = 2482ns;

slave_timing[3][128+31].info_corner          = 1;
slave_timing[3][128+31].info_temp__j__       = -40;
slave_timing[3][128+31].info_i__quite_rec__  = 0.040000000;
slave_timing[3][128+31].info_dtr__ib__       = 1;
slave_timing[3][128+31].info_i__offset_rec__ = 0.000000000;
slave_timing[3][128+31].info_i__max_slave__  = 0.025000000;
slave_timing[3][128+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][128+31].info_r__dsi_bus__    = 5.000;

slave_timing[3][128+31].t_rxd1[0][1] = 2703ns;
slave_timing[3][128+31].t_rxd1[1][0] = 2758ns;
slave_timing[3][128+31].t_rxd1[0][2] = 2036ns;
slave_timing[3][128+31].t_rxd1[2][0] = 3345ns;
slave_timing[3][128+31].t_rxd2[0][2] = 3240ns;
slave_timing[3][128+31].t_rxd2[2][0] = 2067ns;
slave_timing[3][128+31].t_rxd2[1][2] = 2631ns;
slave_timing[3][128+31].t_rxd2[2][1] = 2762ns;

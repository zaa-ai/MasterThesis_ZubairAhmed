
slave_timing[2][160+0].info_corner          = 2;
slave_timing[2][160+0].info_temp__j__       = -40;
slave_timing[2][160+0].info_i__quite_rec__  = 0.006000000;
slave_timing[2][160+0].info_dtr__ib__       = -1;
slave_timing[2][160+0].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+0].info_i__max_slave__  = 0.023000000;
slave_timing[2][160+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][160+0].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+0].t_rxd1[0][1] = 2192ns;
slave_timing[2][160+0].t_rxd1[1][0] = 2207ns;
slave_timing[2][160+0].t_rxd1[0][2] = 1649ns;
slave_timing[2][160+0].t_rxd1[2][0] = 2687ns;
slave_timing[2][160+0].t_rxd2[0][2] = 2640ns;
slave_timing[2][160+0].t_rxd2[2][0] = 1664ns;
slave_timing[2][160+0].t_rxd2[1][2] = 2174ns;
slave_timing[2][160+0].t_rxd2[2][1] = 2197ns;

slave_timing[2][160+1].info_corner          = 2;
slave_timing[2][160+1].info_temp__j__       = -40;
slave_timing[2][160+1].info_i__quite_rec__  = 0.006000000;
slave_timing[2][160+1].info_dtr__ib__       = -1;
slave_timing[2][160+1].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+1].info_i__max_slave__  = 0.025000000;
slave_timing[2][160+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][160+1].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+1].t_rxd1[0][1] = 2110ns;
slave_timing[2][160+1].t_rxd1[1][0] = 2276ns;
slave_timing[2][160+1].t_rxd1[0][2] = 1604ns;
slave_timing[2][160+1].t_rxd1[2][0] = 2732ns;
slave_timing[2][160+1].t_rxd2[0][2] = 2497ns;
slave_timing[2][160+1].t_rxd2[2][0] = 1780ns;
slave_timing[2][160+1].t_rxd2[1][2] = 1941ns;
slave_timing[2][160+1].t_rxd2[2][1] = 2417ns;

slave_timing[2][160+2].info_corner          = 2;
slave_timing[2][160+2].info_temp__j__       = -40;
slave_timing[2][160+2].info_i__quite_rec__  = 0.006000000;
slave_timing[2][160+2].info_dtr__ib__       = 1;
slave_timing[2][160+2].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+2].info_i__max_slave__  = 0.023000000;
slave_timing[2][160+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][160+2].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+2].t_rxd1[0][1] = 2258ns;
slave_timing[2][160+2].t_rxd1[1][0] = 2159ns;
slave_timing[2][160+2].t_rxd1[0][2] = 1684ns;
slave_timing[2][160+2].t_rxd1[2][0] = 2653ns;
slave_timing[2][160+2].t_rxd2[0][2] = 2778ns;
slave_timing[2][160+2].t_rxd2[2][0] = 1563ns;
slave_timing[2][160+2].t_rxd2[1][2] = 2366ns;
slave_timing[2][160+2].t_rxd2[2][1] = 2021ns;

slave_timing[2][160+3].info_corner          = 2;
slave_timing[2][160+3].info_temp__j__       = -40;
slave_timing[2][160+3].info_i__quite_rec__  = 0.006000000;
slave_timing[2][160+3].info_dtr__ib__       = 1;
slave_timing[2][160+3].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+3].info_i__max_slave__  = 0.025000000;
slave_timing[2][160+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][160+3].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+3].t_rxd1[0][1] = 2165ns;
slave_timing[2][160+3].t_rxd1[1][0] = 2228ns;
slave_timing[2][160+3].t_rxd1[0][2] = 1640ns;
slave_timing[2][160+3].t_rxd1[2][0] = 2697ns;
slave_timing[2][160+3].t_rxd2[0][2] = 2601ns;
slave_timing[2][160+3].t_rxd2[2][0] = 1696ns;
slave_timing[2][160+3].t_rxd2[1][2] = 2134ns;
slave_timing[2][160+3].t_rxd2[2][1] = 2217ns;

slave_timing[2][160+4].info_corner          = 2;
slave_timing[2][160+4].info_temp__j__       = -40;
slave_timing[2][160+4].info_i__quite_rec__  = 0.006000000;
slave_timing[2][160+4].info_dtr__ib__       = -1;
slave_timing[2][160+4].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+4].info_i__max_slave__  = 0.023000000;
slave_timing[2][160+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][160+4].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+4].t_rxd1[0][1] = 2263ns;
slave_timing[2][160+4].t_rxd1[1][0] = 2277ns;
slave_timing[2][160+4].t_rxd1[0][2] = 1703ns;
slave_timing[2][160+4].t_rxd1[2][0] = 2752ns;
slave_timing[2][160+4].t_rxd2[0][2] = 2654ns;
slave_timing[2][160+4].t_rxd2[2][0] = 1673ns;
slave_timing[2][160+4].t_rxd2[1][2] = 2182ns;
slave_timing[2][160+4].t_rxd2[2][1] = 2203ns;

slave_timing[2][160+5].info_corner          = 2;
slave_timing[2][160+5].info_temp__j__       = -40;
slave_timing[2][160+5].info_i__quite_rec__  = 0.006000000;
slave_timing[2][160+5].info_dtr__ib__       = -1;
slave_timing[2][160+5].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+5].info_i__max_slave__  = 0.025000000;
slave_timing[2][160+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][160+5].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+5].t_rxd1[0][1] = 2184ns;
slave_timing[2][160+5].t_rxd1[1][0] = 2351ns;
slave_timing[2][160+5].t_rxd1[0][2] = 1667ns;
slave_timing[2][160+5].t_rxd1[2][0] = 2792ns;
slave_timing[2][160+5].t_rxd2[0][2] = 2512ns;
slave_timing[2][160+5].t_rxd2[2][0] = 1793ns;
slave_timing[2][160+5].t_rxd2[1][2] = 1957ns;
slave_timing[2][160+5].t_rxd2[2][1] = 2437ns;

slave_timing[2][160+6].info_corner          = 2;
slave_timing[2][160+6].info_temp__j__       = -40;
slave_timing[2][160+6].info_i__quite_rec__  = 0.006000000;
slave_timing[2][160+6].info_dtr__ib__       = 1;
slave_timing[2][160+6].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+6].info_i__max_slave__  = 0.023000000;
slave_timing[2][160+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][160+6].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+6].t_rxd1[0][1] = 2311ns;
slave_timing[2][160+6].t_rxd1[1][0] = 2223ns;
slave_timing[2][160+6].t_rxd1[0][2] = 1742ns;
slave_timing[2][160+6].t_rxd1[2][0] = 2714ns;
slave_timing[2][160+6].t_rxd2[0][2] = 2788ns;
slave_timing[2][160+6].t_rxd2[2][0] = 1577ns;
slave_timing[2][160+6].t_rxd2[1][2] = 2375ns;
slave_timing[2][160+6].t_rxd2[2][1] = 1997ns;

slave_timing[2][160+7].info_corner          = 2;
slave_timing[2][160+7].info_temp__j__       = -40;
slave_timing[2][160+7].info_i__quite_rec__  = 0.006000000;
slave_timing[2][160+7].info_dtr__ib__       = 1;
slave_timing[2][160+7].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+7].info_i__max_slave__  = 0.025000000;
slave_timing[2][160+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][160+7].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+7].t_rxd1[0][1] = 2219ns;
slave_timing[2][160+7].t_rxd1[1][0] = 2291ns;
slave_timing[2][160+7].t_rxd1[0][2] = 1691ns;
slave_timing[2][160+7].t_rxd1[2][0] = 2757ns;
slave_timing[2][160+7].t_rxd2[0][2] = 2612ns;
slave_timing[2][160+7].t_rxd2[2][0] = 1705ns;
slave_timing[2][160+7].t_rxd2[1][2] = 2114ns;
slave_timing[2][160+7].t_rxd2[2][1] = 2265ns;

slave_timing[2][160+8].info_corner          = 2;
slave_timing[2][160+8].info_temp__j__       = -40;
slave_timing[2][160+8].info_i__quite_rec__  = 0.003000000;
slave_timing[2][160+8].info_dtr__ib__       = -1;
slave_timing[2][160+8].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+8].info_i__max_slave__  = 0.023000000;
slave_timing[2][160+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][160+8].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+8].t_rxd1[0][1] = 2173ns;
slave_timing[2][160+8].t_rxd1[1][0] = 2217ns;
slave_timing[2][160+8].t_rxd1[0][2] = 1645ns;
slave_timing[2][160+8].t_rxd1[2][0] = 2691ns;
slave_timing[2][160+8].t_rxd2[0][2] = 2637ns;
slave_timing[2][160+8].t_rxd2[2][0] = 1669ns;
slave_timing[2][160+8].t_rxd2[1][2] = 2180ns;
slave_timing[2][160+8].t_rxd2[2][1] = 2183ns;

slave_timing[2][160+9].info_corner          = 2;
slave_timing[2][160+9].info_temp__j__       = -40;
slave_timing[2][160+9].info_i__quite_rec__  = 0.003000000;
slave_timing[2][160+9].info_dtr__ib__       = -1;
slave_timing[2][160+9].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+9].info_i__max_slave__  = 0.025000000;
slave_timing[2][160+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][160+9].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+9].t_rxd1[0][1] = 2098ns;
slave_timing[2][160+9].t_rxd1[1][0] = 2279ns;
slave_timing[2][160+9].t_rxd1[0][2] = 1596ns;
slave_timing[2][160+9].t_rxd1[2][0] = 2739ns;
slave_timing[2][160+9].t_rxd2[0][2] = 2492ns;
slave_timing[2][160+9].t_rxd2[2][0] = 1786ns;
slave_timing[2][160+9].t_rxd2[1][2] = 1926ns;
slave_timing[2][160+9].t_rxd2[2][1] = 2442ns;

slave_timing[2][160+10].info_corner          = 2;
slave_timing[2][160+10].info_temp__j__       = -40;
slave_timing[2][160+10].info_i__quite_rec__  = 0.003000000;
slave_timing[2][160+10].info_dtr__ib__       = 1;
slave_timing[2][160+10].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+10].info_i__max_slave__  = 0.023000000;
slave_timing[2][160+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][160+10].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+10].t_rxd1[0][1] = 2238ns;
slave_timing[2][160+10].t_rxd1[1][0] = 2162ns;
slave_timing[2][160+10].t_rxd1[0][2] = 1678ns;
slave_timing[2][160+10].t_rxd1[2][0] = 2655ns;
slave_timing[2][160+10].t_rxd2[0][2] = 2767ns;
slave_timing[2][160+10].t_rxd2[2][0] = 1565ns;
slave_timing[2][160+10].t_rxd2[1][2] = 2352ns;
slave_timing[2][160+10].t_rxd2[2][1] = 2035ns;

slave_timing[2][160+11].info_corner          = 2;
slave_timing[2][160+11].info_temp__j__       = -40;
slave_timing[2][160+11].info_i__quite_rec__  = 0.003000000;
slave_timing[2][160+11].info_dtr__ib__       = 1;
slave_timing[2][160+11].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+11].info_i__max_slave__  = 0.025000000;
slave_timing[2][160+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][160+11].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+11].t_rxd1[0][1] = 2156ns;
slave_timing[2][160+11].t_rxd1[1][0] = 2236ns;
slave_timing[2][160+11].t_rxd1[0][2] = 1629ns;
slave_timing[2][160+11].t_rxd1[2][0] = 2702ns;
slave_timing[2][160+11].t_rxd2[0][2] = 2594ns;
slave_timing[2][160+11].t_rxd2[2][0] = 1704ns;
slave_timing[2][160+11].t_rxd2[1][2] = 2094ns;
slave_timing[2][160+11].t_rxd2[2][1] = 2279ns;

slave_timing[2][160+12].info_corner          = 2;
slave_timing[2][160+12].info_temp__j__       = -40;
slave_timing[2][160+12].info_i__quite_rec__  = 0.003000000;
slave_timing[2][160+12].info_dtr__ib__       = -1;
slave_timing[2][160+12].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+12].info_i__max_slave__  = 0.023000000;
slave_timing[2][160+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][160+12].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+12].t_rxd1[0][1] = 2240ns;
slave_timing[2][160+12].t_rxd1[1][0] = 2290ns;
slave_timing[2][160+12].t_rxd1[0][2] = 1704ns;
slave_timing[2][160+12].t_rxd1[2][0] = 2757ns;
slave_timing[2][160+12].t_rxd2[0][2] = 2649ns;
slave_timing[2][160+12].t_rxd2[2][0] = 1687ns;
slave_timing[2][160+12].t_rxd2[1][2] = 2193ns;
slave_timing[2][160+12].t_rxd2[2][1] = 2192ns;

slave_timing[2][160+13].info_corner          = 2;
slave_timing[2][160+13].info_temp__j__       = -40;
slave_timing[2][160+13].info_i__quite_rec__  = 0.003000000;
slave_timing[2][160+13].info_dtr__ib__       = -1;
slave_timing[2][160+13].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+13].info_i__max_slave__  = 0.025000000;
slave_timing[2][160+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][160+13].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+13].t_rxd1[0][1] = 2166ns;
slave_timing[2][160+13].t_rxd1[1][0] = 2361ns;
slave_timing[2][160+13].t_rxd1[0][2] = 1661ns;
slave_timing[2][160+13].t_rxd1[2][0] = 2800ns;
slave_timing[2][160+13].t_rxd2[0][2] = 2506ns;
slave_timing[2][160+13].t_rxd2[2][0] = 1799ns;
slave_timing[2][160+13].t_rxd2[1][2] = 1932ns;
slave_timing[2][160+13].t_rxd2[2][1] = 2456ns;

slave_timing[2][160+14].info_corner          = 2;
slave_timing[2][160+14].info_temp__j__       = -40;
slave_timing[2][160+14].info_i__quite_rec__  = 0.003000000;
slave_timing[2][160+14].info_dtr__ib__       = 1;
slave_timing[2][160+14].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+14].info_i__max_slave__  = 0.023000000;
slave_timing[2][160+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][160+14].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+14].t_rxd1[0][1] = 2297ns;
slave_timing[2][160+14].t_rxd1[1][0] = 2216ns;
slave_timing[2][160+14].t_rxd1[0][2] = 1729ns;
slave_timing[2][160+14].t_rxd1[2][0] = 2718ns;
slave_timing[2][160+14].t_rxd2[0][2] = 2780ns;
slave_timing[2][160+14].t_rxd2[2][0] = 1585ns;
slave_timing[2][160+14].t_rxd2[1][2] = 2360ns;
slave_timing[2][160+14].t_rxd2[2][1] = 2047ns;

slave_timing[2][160+15].info_corner          = 2;
slave_timing[2][160+15].info_temp__j__       = -40;
slave_timing[2][160+15].info_i__quite_rec__  = 0.003000000;
slave_timing[2][160+15].info_dtr__ib__       = 1;
slave_timing[2][160+15].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+15].info_i__max_slave__  = 0.025000000;
slave_timing[2][160+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][160+15].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+15].t_rxd1[0][1] = 2216ns;
slave_timing[2][160+15].t_rxd1[1][0] = 2295ns;
slave_timing[2][160+15].t_rxd1[0][2] = 1686ns;
slave_timing[2][160+15].t_rxd1[2][0] = 2764ns;
slave_timing[2][160+15].t_rxd2[0][2] = 2605ns;
slave_timing[2][160+15].t_rxd2[2][0] = 1717ns;
slave_timing[2][160+15].t_rxd2[1][2] = 2104ns;
slave_timing[2][160+15].t_rxd2[2][1] = 2263ns;

slave_timing[2][160+16].info_corner          = 2;
slave_timing[2][160+16].info_temp__j__       = -40;
slave_timing[2][160+16].info_i__quite_rec__  = 0.000000000;
slave_timing[2][160+16].info_dtr__ib__       = -1;
slave_timing[2][160+16].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+16].info_i__max_slave__  = 0.023000000;
slave_timing[2][160+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][160+16].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+16].t_rxd1[0][1] = 2186ns;
slave_timing[2][160+16].t_rxd1[1][0] = 2205ns;
slave_timing[2][160+16].t_rxd1[0][2] = 1656ns;
slave_timing[2][160+16].t_rxd1[2][0] = 2681ns;
slave_timing[2][160+16].t_rxd2[0][2] = 2646ns;
slave_timing[2][160+16].t_rxd2[2][0] = 1657ns;
slave_timing[2][160+16].t_rxd2[1][2] = 2156ns;
slave_timing[2][160+16].t_rxd2[2][1] = 2198ns;

slave_timing[2][160+17].info_corner          = 2;
slave_timing[2][160+17].info_temp__j__       = -40;
slave_timing[2][160+17].info_i__quite_rec__  = 0.000000000;
slave_timing[2][160+17].info_dtr__ib__       = -1;
slave_timing[2][160+17].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+17].info_i__max_slave__  = 0.025000000;
slave_timing[2][160+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][160+17].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+17].t_rxd1[0][1] = 2109ns;
slave_timing[2][160+17].t_rxd1[1][0] = 2267ns;
slave_timing[2][160+17].t_rxd1[0][2] = 1609ns;
slave_timing[2][160+17].t_rxd1[2][0] = 2725ns;
slave_timing[2][160+17].t_rxd2[0][2] = 2500ns;
slave_timing[2][160+17].t_rxd2[2][0] = 1777ns;
slave_timing[2][160+17].t_rxd2[1][2] = 1946ns;
slave_timing[2][160+17].t_rxd2[2][1] = 2428ns;

slave_timing[2][160+18].info_corner          = 2;
slave_timing[2][160+18].info_temp__j__       = -40;
slave_timing[2][160+18].info_i__quite_rec__  = 0.000000000;
slave_timing[2][160+18].info_dtr__ib__       = 1;
slave_timing[2][160+18].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+18].info_i__max_slave__  = 0.023000000;
slave_timing[2][160+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][160+18].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+18].t_rxd1[0][1] = 2261ns;
slave_timing[2][160+18].t_rxd1[1][0] = 2147ns;
slave_timing[2][160+18].t_rxd1[0][2] = 1692ns;
slave_timing[2][160+18].t_rxd1[2][0] = 2640ns;
slave_timing[2][160+18].t_rxd2[0][2] = 2778ns;
slave_timing[2][160+18].t_rxd2[2][0] = 1555ns;
slave_timing[2][160+18].t_rxd2[1][2] = 2368ns;
slave_timing[2][160+18].t_rxd2[2][1] = 2006ns;

slave_timing[2][160+19].info_corner          = 2;
slave_timing[2][160+19].info_temp__j__       = -40;
slave_timing[2][160+19].info_i__quite_rec__  = 0.000000000;
slave_timing[2][160+19].info_dtr__ib__       = 1;
slave_timing[2][160+19].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+19].info_i__max_slave__  = 0.025000000;
slave_timing[2][160+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][160+19].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+19].t_rxd1[0][1] = 2166ns;
slave_timing[2][160+19].t_rxd1[1][0] = 2214ns;
slave_timing[2][160+19].t_rxd1[0][2] = 1641ns;
slave_timing[2][160+19].t_rxd1[2][0] = 2694ns;
slave_timing[2][160+19].t_rxd2[0][2] = 2603ns;
slave_timing[2][160+19].t_rxd2[2][0] = 1690ns;
slave_timing[2][160+19].t_rxd2[1][2] = 2110ns;
slave_timing[2][160+19].t_rxd2[2][1] = 2246ns;

slave_timing[2][160+20].info_corner          = 2;
slave_timing[2][160+20].info_temp__j__       = -40;
slave_timing[2][160+20].info_i__quite_rec__  = 0.000000000;
slave_timing[2][160+20].info_dtr__ib__       = -1;
slave_timing[2][160+20].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+20].info_i__max_slave__  = 0.023000000;
slave_timing[2][160+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][160+20].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+20].t_rxd1[0][1] = 2262ns;
slave_timing[2][160+20].t_rxd1[1][0] = 2262ns;
slave_timing[2][160+20].t_rxd1[0][2] = 1720ns;
slave_timing[2][160+20].t_rxd1[2][0] = 2747ns;
slave_timing[2][160+20].t_rxd2[0][2] = 2658ns;
slave_timing[2][160+20].t_rxd2[2][0] = 1677ns;
slave_timing[2][160+20].t_rxd2[1][2] = 2180ns;
slave_timing[2][160+20].t_rxd2[2][1] = 2200ns;

slave_timing[2][160+21].info_corner          = 2;
slave_timing[2][160+21].info_temp__j__       = -40;
slave_timing[2][160+21].info_i__quite_rec__  = 0.000000000;
slave_timing[2][160+21].info_dtr__ib__       = -1;
slave_timing[2][160+21].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+21].info_i__max_slave__  = 0.025000000;
slave_timing[2][160+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][160+21].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+21].t_rxd1[0][1] = 2179ns;
slave_timing[2][160+21].t_rxd1[1][0] = 2333ns;
slave_timing[2][160+21].t_rxd1[0][2] = 1672ns;
slave_timing[2][160+21].t_rxd1[2][0] = 2792ns;
slave_timing[2][160+21].t_rxd2[0][2] = 2514ns;
slave_timing[2][160+21].t_rxd2[2][0] = 1791ns;
slave_timing[2][160+21].t_rxd2[1][2] = 1964ns;
slave_timing[2][160+21].t_rxd2[2][1] = 2438ns;

slave_timing[2][160+22].info_corner          = 2;
slave_timing[2][160+22].info_temp__j__       = -40;
slave_timing[2][160+22].info_i__quite_rec__  = 0.000000000;
slave_timing[2][160+22].info_dtr__ib__       = 1;
slave_timing[2][160+22].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+22].info_i__max_slave__  = 0.023000000;
slave_timing[2][160+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][160+22].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+22].t_rxd1[0][1] = 2328ns;
slave_timing[2][160+22].t_rxd1[1][0] = 2205ns;
slave_timing[2][160+22].t_rxd1[0][2] = 1746ns;
slave_timing[2][160+22].t_rxd1[2][0] = 2705ns;
slave_timing[2][160+22].t_rxd2[0][2] = 2788ns;
slave_timing[2][160+22].t_rxd2[2][0] = 1565ns;
slave_timing[2][160+22].t_rxd2[1][2] = 2404ns;
slave_timing[2][160+22].t_rxd2[2][1] = 1988ns;

slave_timing[2][160+23].info_corner          = 2;
slave_timing[2][160+23].info_temp__j__       = -40;
slave_timing[2][160+23].info_i__quite_rec__  = 0.000000000;
slave_timing[2][160+23].info_dtr__ib__       = 1;
slave_timing[2][160+23].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+23].info_i__max_slave__  = 0.025000000;
slave_timing[2][160+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][160+23].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+23].t_rxd1[0][1] = 2228ns;
slave_timing[2][160+23].t_rxd1[1][0] = 2277ns;
slave_timing[2][160+23].t_rxd1[0][2] = 1700ns;
slave_timing[2][160+23].t_rxd1[2][0] = 2751ns;
slave_timing[2][160+23].t_rxd2[0][2] = 2619ns;
slave_timing[2][160+23].t_rxd2[2][0] = 1697ns;
slave_timing[2][160+23].t_rxd2[1][2] = 2128ns;
slave_timing[2][160+23].t_rxd2[2][1] = 2218ns;

slave_timing[2][160+24].info_corner          = 2;
slave_timing[2][160+24].info_temp__j__       = -40;
slave_timing[2][160+24].info_i__quite_rec__  = 0.040000000;
slave_timing[2][160+24].info_dtr__ib__       = -1;
slave_timing[2][160+24].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+24].info_i__max_slave__  = 0.023000000;
slave_timing[2][160+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][160+24].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+24].t_rxd1[0][1] = 2192ns;
slave_timing[2][160+24].t_rxd1[1][0] = 2188ns;
slave_timing[2][160+24].t_rxd1[0][2] = 1650ns;
slave_timing[2][160+24].t_rxd1[2][0] = 2672ns;
slave_timing[2][160+24].t_rxd2[0][2] = 2644ns;
slave_timing[2][160+24].t_rxd2[2][0] = 1654ns;
slave_timing[2][160+24].t_rxd2[1][2] = 2166ns;
slave_timing[2][160+24].t_rxd2[2][1] = 2189ns;

slave_timing[2][160+25].info_corner          = 2;
slave_timing[2][160+25].info_temp__j__       = -40;
slave_timing[2][160+25].info_i__quite_rec__  = 0.040000000;
slave_timing[2][160+25].info_dtr__ib__       = -1;
slave_timing[2][160+25].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+25].info_i__max_slave__  = 0.025000000;
slave_timing[2][160+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][160+25].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+25].t_rxd1[0][1] = 2110ns;
slave_timing[2][160+25].t_rxd1[1][0] = 2256ns;
slave_timing[2][160+25].t_rxd1[0][2] = 1604ns;
slave_timing[2][160+25].t_rxd1[2][0] = 2719ns;
slave_timing[2][160+25].t_rxd2[0][2] = 2499ns;
slave_timing[2][160+25].t_rxd2[2][0] = 1775ns;
slave_timing[2][160+25].t_rxd2[1][2] = 1944ns;
slave_timing[2][160+25].t_rxd2[2][1] = 2427ns;

slave_timing[2][160+26].info_corner          = 2;
slave_timing[2][160+26].info_temp__j__       = -40;
slave_timing[2][160+26].info_i__quite_rec__  = 0.040000000;
slave_timing[2][160+26].info_dtr__ib__       = 1;
slave_timing[2][160+26].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+26].info_i__max_slave__  = 0.023000000;
slave_timing[2][160+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][160+26].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+26].t_rxd1[0][1] = 2240ns;
slave_timing[2][160+26].t_rxd1[1][0] = 2153ns;
slave_timing[2][160+26].t_rxd1[0][2] = 1681ns;
slave_timing[2][160+26].t_rxd1[2][0] = 2645ns;
slave_timing[2][160+26].t_rxd2[0][2] = 2766ns;
slave_timing[2][160+26].t_rxd2[2][0] = 1555ns;
slave_timing[2][160+26].t_rxd2[1][2] = 2358ns;
slave_timing[2][160+26].t_rxd2[2][1] = 2026ns;

slave_timing[2][160+27].info_corner          = 2;
slave_timing[2][160+27].info_temp__j__       = -40;
slave_timing[2][160+27].info_i__quite_rec__  = 0.040000000;
slave_timing[2][160+27].info_dtr__ib__       = 1;
slave_timing[2][160+27].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+27].info_i__max_slave__  = 0.025000000;
slave_timing[2][160+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][160+27].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+27].t_rxd1[0][1] = 2160ns;
slave_timing[2][160+27].t_rxd1[1][0] = 2217ns;
slave_timing[2][160+27].t_rxd1[0][2] = 1632ns;
slave_timing[2][160+27].t_rxd1[2][0] = 2697ns;
slave_timing[2][160+27].t_rxd2[0][2] = 2601ns;
slave_timing[2][160+27].t_rxd2[2][0] = 1697ns;
slave_timing[2][160+27].t_rxd2[1][2] = 2103ns;
slave_timing[2][160+27].t_rxd2[2][1] = 2255ns;

slave_timing[2][160+28].info_corner          = 2;
slave_timing[2][160+28].info_temp__j__       = -40;
slave_timing[2][160+28].info_i__quite_rec__  = 0.040000000;
slave_timing[2][160+28].info_dtr__ib__       = -1;
slave_timing[2][160+28].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+28].info_i__max_slave__  = 0.023000000;
slave_timing[2][160+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][160+28].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+28].t_rxd1[0][1] = 2226ns;
slave_timing[2][160+28].t_rxd1[1][0] = 2229ns;
slave_timing[2][160+28].t_rxd1[0][2] = 1688ns;
slave_timing[2][160+28].t_rxd1[2][0] = 2712ns;
slave_timing[2][160+28].t_rxd2[0][2] = 2667ns;
slave_timing[2][160+28].t_rxd2[2][0] = 1674ns;
slave_timing[2][160+28].t_rxd2[1][2] = 2186ns;
slave_timing[2][160+28].t_rxd2[2][1] = 2202ns;

slave_timing[2][160+29].info_corner          = 2;
slave_timing[2][160+29].info_temp__j__       = -40;
slave_timing[2][160+29].info_i__quite_rec__  = 0.040000000;
slave_timing[2][160+29].info_dtr__ib__       = -1;
slave_timing[2][160+29].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+29].info_i__max_slave__  = 0.025000000;
slave_timing[2][160+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][160+29].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+29].t_rxd1[0][1] = 2133ns;
slave_timing[2][160+29].t_rxd1[1][0] = 2306ns;
slave_timing[2][160+29].t_rxd1[0][2] = 1640ns;
slave_timing[2][160+29].t_rxd1[2][0] = 2758ns;
slave_timing[2][160+29].t_rxd2[0][2] = 2511ns;
slave_timing[2][160+29].t_rxd2[2][0] = 1788ns;
slave_timing[2][160+29].t_rxd2[1][2] = 1953ns;
slave_timing[2][160+29].t_rxd2[2][1] = 2433ns;

slave_timing[2][160+30].info_corner          = 2;
slave_timing[2][160+30].info_temp__j__       = -40;
slave_timing[2][160+30].info_i__quite_rec__  = 0.040000000;
slave_timing[2][160+30].info_dtr__ib__       = 1;
slave_timing[2][160+30].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+30].info_i__max_slave__  = 0.023000000;
slave_timing[2][160+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][160+30].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+30].t_rxd1[0][1] = 2276ns;
slave_timing[2][160+30].t_rxd1[1][0] = 2196ns;
slave_timing[2][160+30].t_rxd1[0][2] = 1704ns;
slave_timing[2][160+30].t_rxd1[2][0] = 2684ns;
slave_timing[2][160+30].t_rxd2[0][2] = 2785ns;
slave_timing[2][160+30].t_rxd2[2][0] = 1576ns;
slave_timing[2][160+30].t_rxd2[1][2] = 2369ns;
slave_timing[2][160+30].t_rxd2[2][1] = 2034ns;

slave_timing[2][160+31].info_corner          = 2;
slave_timing[2][160+31].info_temp__j__       = -40;
slave_timing[2][160+31].info_i__quite_rec__  = 0.040000000;
slave_timing[2][160+31].info_dtr__ib__       = 1;
slave_timing[2][160+31].info_i__offset_rec__ = 0.000000000;
slave_timing[2][160+31].info_i__max_slave__  = 0.025000000;
slave_timing[2][160+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][160+31].info_r__dsi_bus__    = 5.000;

slave_timing[2][160+31].t_rxd1[0][1] = 2190ns;
slave_timing[2][160+31].t_rxd1[1][0] = 2265ns;
slave_timing[2][160+31].t_rxd1[0][2] = 1662ns;
slave_timing[2][160+31].t_rxd1[2][0] = 2728ns;
slave_timing[2][160+31].t_rxd2[0][2] = 2612ns;
slave_timing[2][160+31].t_rxd2[2][0] = 1708ns;
slave_timing[2][160+31].t_rxd2[1][2] = 2113ns;
slave_timing[2][160+31].t_rxd2[2][1] = 2263ns;


slave_timing[3][160+0].info_corner          = 2;
slave_timing[3][160+0].info_temp__j__       = -40;
slave_timing[3][160+0].info_i__quite_rec__  = 0.006000000;
slave_timing[3][160+0].info_dtr__ib__       = -1;
slave_timing[3][160+0].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+0].info_i__max_slave__  = 0.023000000;
slave_timing[3][160+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][160+0].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+0].t_rxd1[0][1] = 2737ns;
slave_timing[3][160+0].t_rxd1[1][0] = 2740ns;
slave_timing[3][160+0].t_rxd1[0][2] = 2047ns;
slave_timing[3][160+0].t_rxd1[2][0] = 3342ns;
slave_timing[3][160+0].t_rxd2[0][2] = 3313ns;
slave_timing[3][160+0].t_rxd2[2][0] = 2050ns;
slave_timing[3][160+0].t_rxd2[1][2] = 2720ns;
slave_timing[3][160+0].t_rxd2[2][1] = 2729ns;

slave_timing[3][160+1].info_corner          = 2;
slave_timing[3][160+1].info_temp__j__       = -40;
slave_timing[3][160+1].info_i__quite_rec__  = 0.006000000;
slave_timing[3][160+1].info_dtr__ib__       = -1;
slave_timing[3][160+1].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+1].info_i__max_slave__  = 0.025000000;
slave_timing[3][160+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][160+1].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+1].t_rxd1[0][1] = 2633ns;
slave_timing[3][160+1].t_rxd1[1][0] = 2823ns;
slave_timing[3][160+1].t_rxd1[0][2] = 1986ns;
slave_timing[3][160+1].t_rxd1[2][0] = 3397ns;
slave_timing[3][160+1].t_rxd2[0][2] = 3124ns;
slave_timing[3][160+1].t_rxd2[2][0] = 2197ns;
slave_timing[3][160+1].t_rxd2[1][2] = 2430ns;
slave_timing[3][160+1].t_rxd2[2][1] = 2976ns;

slave_timing[3][160+2].info_corner          = 2;
slave_timing[3][160+2].info_temp__j__       = -40;
slave_timing[3][160+2].info_i__quite_rec__  = 0.006000000;
slave_timing[3][160+2].info_dtr__ib__       = 1;
slave_timing[3][160+2].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+2].info_i__max_slave__  = 0.023000000;
slave_timing[3][160+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][160+2].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+2].t_rxd1[0][1] = 2823ns;
slave_timing[3][160+2].t_rxd1[1][0] = 2678ns;
slave_timing[3][160+2].t_rxd1[0][2] = 2096ns;
slave_timing[3][160+2].t_rxd1[2][0] = 3302ns;
slave_timing[3][160+2].t_rxd2[0][2] = 3484ns;
slave_timing[3][160+2].t_rxd2[2][0] = 1919ns;
slave_timing[3][160+2].t_rxd2[1][2] = 2968ns;
slave_timing[3][160+2].t_rxd2[2][1] = 2475ns;

slave_timing[3][160+3].info_corner          = 2;
slave_timing[3][160+3].info_temp__j__       = -40;
slave_timing[3][160+3].info_i__quite_rec__  = 0.006000000;
slave_timing[3][160+3].info_dtr__ib__       = 1;
slave_timing[3][160+3].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+3].info_i__max_slave__  = 0.025000000;
slave_timing[3][160+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][160+3].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+3].t_rxd1[0][1] = 2709ns;
slave_timing[3][160+3].t_rxd1[1][0] = 2762ns;
slave_timing[3][160+3].t_rxd1[0][2] = 2028ns;
slave_timing[3][160+3].t_rxd1[2][0] = 3354ns;
slave_timing[3][160+3].t_rxd2[0][2] = 3253ns;
slave_timing[3][160+3].t_rxd2[2][0] = 2090ns;
slave_timing[3][160+3].t_rxd2[1][2] = 2676ns;
slave_timing[3][160+3].t_rxd2[2][1] = 2763ns;

slave_timing[3][160+4].info_corner          = 2;
slave_timing[3][160+4].info_temp__j__       = -40;
slave_timing[3][160+4].info_i__quite_rec__  = 0.006000000;
slave_timing[3][160+4].info_dtr__ib__       = -1;
slave_timing[3][160+4].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+4].info_i__max_slave__  = 0.023000000;
slave_timing[3][160+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][160+4].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+4].t_rxd1[0][1] = 2809ns;
slave_timing[3][160+4].t_rxd1[1][0] = 2808ns;
slave_timing[3][160+4].t_rxd1[0][2] = 2110ns;
slave_timing[3][160+4].t_rxd1[2][0] = 3405ns;
slave_timing[3][160+4].t_rxd2[0][2] = 3323ns;
slave_timing[3][160+4].t_rxd2[2][0] = 2058ns;
slave_timing[3][160+4].t_rxd2[1][2] = 2731ns;
slave_timing[3][160+4].t_rxd2[2][1] = 2741ns;

slave_timing[3][160+5].info_corner          = 2;
slave_timing[3][160+5].info_temp__j__       = -40;
slave_timing[3][160+5].info_i__quite_rec__  = 0.006000000;
slave_timing[3][160+5].info_dtr__ib__       = -1;
slave_timing[3][160+5].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+5].info_i__max_slave__  = 0.025000000;
slave_timing[3][160+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][160+5].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+5].t_rxd1[0][1] = 2692ns;
slave_timing[3][160+5].t_rxd1[1][0] = 2891ns;
slave_timing[3][160+5].t_rxd1[0][2] = 2045ns;
slave_timing[3][160+5].t_rxd1[2][0] = 3460ns;
slave_timing[3][160+5].t_rxd2[0][2] = 3135ns;
slave_timing[3][160+5].t_rxd2[2][0] = 2207ns;
slave_timing[3][160+5].t_rxd2[1][2] = 2442ns;
slave_timing[3][160+5].t_rxd2[2][1] = 3027ns;

slave_timing[3][160+6].info_corner          = 2;
slave_timing[3][160+6].info_temp__j__       = -40;
slave_timing[3][160+6].info_i__quite_rec__  = 0.006000000;
slave_timing[3][160+6].info_dtr__ib__       = 1;
slave_timing[3][160+6].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+6].info_i__max_slave__  = 0.023000000;
slave_timing[3][160+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][160+6].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+6].t_rxd1[0][1] = 2886ns;
slave_timing[3][160+6].t_rxd1[1][0] = 2739ns;
slave_timing[3][160+6].t_rxd1[0][2] = 2152ns;
slave_timing[3][160+6].t_rxd1[2][0] = 3360ns;
slave_timing[3][160+6].t_rxd2[0][2] = 3494ns;
slave_timing[3][160+6].t_rxd2[2][0] = 1929ns;
slave_timing[3][160+6].t_rxd2[1][2] = 3024ns;
slave_timing[3][160+6].t_rxd2[2][1] = 2485ns;

slave_timing[3][160+7].info_corner          = 2;
slave_timing[3][160+7].info_temp__j__       = -40;
slave_timing[3][160+7].info_i__quite_rec__  = 0.006000000;
slave_timing[3][160+7].info_dtr__ib__       = 1;
slave_timing[3][160+7].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+7].info_i__max_slave__  = 0.025000000;
slave_timing[3][160+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][160+7].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+7].t_rxd1[0][1] = 2769ns;
slave_timing[3][160+7].t_rxd1[1][0] = 2823ns;
slave_timing[3][160+7].t_rxd1[0][2] = 2084ns;
slave_timing[3][160+7].t_rxd1[2][0] = 3418ns;
slave_timing[3][160+7].t_rxd2[0][2] = 3269ns;
slave_timing[3][160+7].t_rxd2[2][0] = 2091ns;
slave_timing[3][160+7].t_rxd2[1][2] = 2648ns;
slave_timing[3][160+7].t_rxd2[2][1] = 2812ns;

slave_timing[3][160+8].info_corner          = 2;
slave_timing[3][160+8].info_temp__j__       = -40;
slave_timing[3][160+8].info_i__quite_rec__  = 0.003000000;
slave_timing[3][160+8].info_dtr__ib__       = -1;
slave_timing[3][160+8].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+8].info_i__max_slave__  = 0.023000000;
slave_timing[3][160+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][160+8].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+8].t_rxd1[0][1] = 2719ns;
slave_timing[3][160+8].t_rxd1[1][0] = 2749ns;
slave_timing[3][160+8].t_rxd1[0][2] = 2037ns;
slave_timing[3][160+8].t_rxd1[2][0] = 3347ns;
slave_timing[3][160+8].t_rxd2[0][2] = 3303ns;
slave_timing[3][160+8].t_rxd2[2][0] = 2060ns;
slave_timing[3][160+8].t_rxd2[1][2] = 2739ns;
slave_timing[3][160+8].t_rxd2[2][1] = 2709ns;

slave_timing[3][160+9].info_corner          = 2;
slave_timing[3][160+9].info_temp__j__       = -40;
slave_timing[3][160+9].info_i__quite_rec__  = 0.003000000;
slave_timing[3][160+9].info_dtr__ib__       = -1;
slave_timing[3][160+9].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+9].info_i__max_slave__  = 0.025000000;
slave_timing[3][160+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][160+9].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+9].t_rxd1[0][1] = 2620ns;
slave_timing[3][160+9].t_rxd1[1][0] = 2833ns;
slave_timing[3][160+9].t_rxd1[0][2] = 1975ns;
slave_timing[3][160+9].t_rxd1[2][0] = 3405ns;
slave_timing[3][160+9].t_rxd2[0][2] = 3107ns;
slave_timing[3][160+9].t_rxd2[2][0] = 2204ns;
slave_timing[3][160+9].t_rxd2[1][2] = 2413ns;
slave_timing[3][160+9].t_rxd2[2][1] = 3038ns;

slave_timing[3][160+10].info_corner          = 2;
slave_timing[3][160+10].info_temp__j__       = -40;
slave_timing[3][160+10].info_i__quite_rec__  = 0.003000000;
slave_timing[3][160+10].info_dtr__ib__       = 1;
slave_timing[3][160+10].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+10].info_i__max_slave__  = 0.023000000;
slave_timing[3][160+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][160+10].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+10].t_rxd1[0][1] = 2807ns;
slave_timing[3][160+10].t_rxd1[1][0] = 2687ns;
slave_timing[3][160+10].t_rxd1[0][2] = 2083ns;
slave_timing[3][160+10].t_rxd1[2][0] = 3306ns;
slave_timing[3][160+10].t_rxd2[0][2] = 3472ns;
slave_timing[3][160+10].t_rxd2[2][0] = 1925ns;
slave_timing[3][160+10].t_rxd2[1][2] = 2950ns;
slave_timing[3][160+10].t_rxd2[2][1] = 2534ns;

slave_timing[3][160+11].info_corner          = 2;
slave_timing[3][160+11].info_temp__j__       = -40;
slave_timing[3][160+11].info_i__quite_rec__  = 0.003000000;
slave_timing[3][160+11].info_dtr__ib__       = 1;
slave_timing[3][160+11].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+11].info_i__max_slave__  = 0.025000000;
slave_timing[3][160+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][160+11].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+11].t_rxd1[0][1] = 2696ns;
slave_timing[3][160+11].t_rxd1[1][0] = 2771ns;
slave_timing[3][160+11].t_rxd1[0][2] = 2014ns;
slave_timing[3][160+11].t_rxd1[2][0] = 3360ns;
slave_timing[3][160+11].t_rxd2[0][2] = 3247ns;
slave_timing[3][160+11].t_rxd2[2][0] = 2098ns;
slave_timing[3][160+11].t_rxd2[1][2] = 2617ns;
slave_timing[3][160+11].t_rxd2[2][1] = 2814ns;

slave_timing[3][160+12].info_corner          = 2;
slave_timing[3][160+12].info_temp__j__       = -40;
slave_timing[3][160+12].info_i__quite_rec__  = 0.003000000;
slave_timing[3][160+12].info_dtr__ib__       = -1;
slave_timing[3][160+12].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+12].info_i__max_slave__  = 0.023000000;
slave_timing[3][160+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][160+12].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+12].t_rxd1[0][1] = 2823ns;
slave_timing[3][160+12].t_rxd1[1][0] = 2781ns;
slave_timing[3][160+12].t_rxd1[0][2] = 2100ns;
slave_timing[3][160+12].t_rxd1[2][0] = 3416ns;
slave_timing[3][160+12].t_rxd2[0][2] = 3309ns;
slave_timing[3][160+12].t_rxd2[2][0] = 2074ns;
slave_timing[3][160+12].t_rxd2[1][2] = 2753ns;
slave_timing[3][160+12].t_rxd2[2][1] = 2718ns;

slave_timing[3][160+13].info_corner          = 2;
slave_timing[3][160+13].info_temp__j__       = -40;
slave_timing[3][160+13].info_i__quite_rec__  = 0.003000000;
slave_timing[3][160+13].info_dtr__ib__       = -1;
slave_timing[3][160+13].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+13].info_i__max_slave__  = 0.025000000;
slave_timing[3][160+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][160+13].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+13].t_rxd1[0][1] = 2684ns;
slave_timing[3][160+13].t_rxd1[1][0] = 2909ns;
slave_timing[3][160+13].t_rxd1[0][2] = 2033ns;
slave_timing[3][160+13].t_rxd1[2][0] = 3470ns;
slave_timing[3][160+13].t_rxd2[0][2] = 3125ns;
slave_timing[3][160+13].t_rxd2[2][0] = 2222ns;
slave_timing[3][160+13].t_rxd2[1][2] = 2427ns;
slave_timing[3][160+13].t_rxd2[2][1] = 3043ns;

slave_timing[3][160+14].info_corner          = 2;
slave_timing[3][160+14].info_temp__j__       = -40;
slave_timing[3][160+14].info_i__quite_rec__  = 0.003000000;
slave_timing[3][160+14].info_dtr__ib__       = 1;
slave_timing[3][160+14].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+14].info_i__max_slave__  = 0.023000000;
slave_timing[3][160+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][160+14].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+14].t_rxd1[0][1] = 2869ns;
slave_timing[3][160+14].t_rxd1[1][0] = 2750ns;
slave_timing[3][160+14].t_rxd1[0][2] = 2141ns;
slave_timing[3][160+14].t_rxd1[2][0] = 3369ns;
slave_timing[3][160+14].t_rxd2[0][2] = 3482ns;
slave_timing[3][160+14].t_rxd2[2][0] = 1940ns;
slave_timing[3][160+14].t_rxd2[1][2] = 2955ns;
slave_timing[3][160+14].t_rxd2[2][1] = 2542ns;

slave_timing[3][160+15].info_corner          = 2;
slave_timing[3][160+15].info_temp__j__       = -40;
slave_timing[3][160+15].info_i__quite_rec__  = 0.003000000;
slave_timing[3][160+15].info_dtr__ib__       = 1;
slave_timing[3][160+15].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+15].info_i__max_slave__  = 0.025000000;
slave_timing[3][160+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][160+15].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+15].t_rxd1[0][1] = 2753ns;
slave_timing[3][160+15].t_rxd1[1][0] = 2835ns;
slave_timing[3][160+15].t_rxd1[0][2] = 2078ns;
slave_timing[3][160+15].t_rxd1[2][0] = 3423ns;
slave_timing[3][160+15].t_rxd2[0][2] = 3259ns;
slave_timing[3][160+15].t_rxd2[2][0] = 2112ns;
slave_timing[3][160+15].t_rxd2[1][2] = 2633ns;
slave_timing[3][160+15].t_rxd2[2][1] = 2830ns;

slave_timing[3][160+16].info_corner          = 2;
slave_timing[3][160+16].info_temp__j__       = -40;
slave_timing[3][160+16].info_i__quite_rec__  = 0.000000000;
slave_timing[3][160+16].info_dtr__ib__       = -1;
slave_timing[3][160+16].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+16].info_i__max_slave__  = 0.023000000;
slave_timing[3][160+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][160+16].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+16].t_rxd1[0][1] = 2744ns;
slave_timing[3][160+16].t_rxd1[1][0] = 2731ns;
slave_timing[3][160+16].t_rxd1[0][2] = 2051ns;
slave_timing[3][160+16].t_rxd1[2][0] = 3335ns;
slave_timing[3][160+16].t_rxd2[0][2] = 3315ns;
slave_timing[3][160+16].t_rxd2[2][0] = 2046ns;
slave_timing[3][160+16].t_rxd2[1][2] = 2730ns;
slave_timing[3][160+16].t_rxd2[2][1] = 2727ns;

slave_timing[3][160+17].info_corner          = 2;
slave_timing[3][160+17].info_temp__j__       = -40;
slave_timing[3][160+17].info_i__quite_rec__  = 0.000000000;
slave_timing[3][160+17].info_dtr__ib__       = -1;
slave_timing[3][160+17].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+17].info_i__max_slave__  = 0.025000000;
slave_timing[3][160+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][160+17].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+17].t_rxd1[0][1] = 2639ns;
slave_timing[3][160+17].t_rxd1[1][0] = 2814ns;
slave_timing[3][160+17].t_rxd1[0][2] = 1983ns;
slave_timing[3][160+17].t_rxd1[2][0] = 3390ns;
slave_timing[3][160+17].t_rxd2[0][2] = 3126ns;
slave_timing[3][160+17].t_rxd2[2][0] = 2194ns;
slave_timing[3][160+17].t_rxd2[1][2] = 2435ns;
slave_timing[3][160+17].t_rxd2[2][1] = 3015ns;

slave_timing[3][160+18].info_corner          = 2;
slave_timing[3][160+18].info_temp__j__       = -40;
slave_timing[3][160+18].info_i__quite_rec__  = 0.000000000;
slave_timing[3][160+18].info_dtr__ib__       = 1;
slave_timing[3][160+18].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+18].info_i__max_slave__  = 0.023000000;
slave_timing[3][160+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][160+18].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+18].t_rxd1[0][1] = 2835ns;
slave_timing[3][160+18].t_rxd1[1][0] = 2663ns;
slave_timing[3][160+18].t_rxd1[0][2] = 2102ns;
slave_timing[3][160+18].t_rxd1[2][0] = 3292ns;
slave_timing[3][160+18].t_rxd2[0][2] = 3494ns;
slave_timing[3][160+18].t_rxd2[2][0] = 1909ns;
slave_timing[3][160+18].t_rxd2[1][2] = 2981ns;
slave_timing[3][160+18].t_rxd2[2][1] = 2495ns;

slave_timing[3][160+19].info_corner          = 2;
slave_timing[3][160+19].info_temp__j__       = -40;
slave_timing[3][160+19].info_i__quite_rec__  = 0.000000000;
slave_timing[3][160+19].info_dtr__ib__       = 1;
slave_timing[3][160+19].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+19].info_i__max_slave__  = 0.025000000;
slave_timing[3][160+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][160+19].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+19].t_rxd1[0][1] = 2718ns;
slave_timing[3][160+19].t_rxd1[1][0] = 2752ns;
slave_timing[3][160+19].t_rxd1[0][2] = 2034ns;
slave_timing[3][160+19].t_rxd1[2][0] = 3348ns;
slave_timing[3][160+19].t_rxd2[0][2] = 3264ns;
slave_timing[3][160+19].t_rxd2[2][0] = 2081ns;
slave_timing[3][160+19].t_rxd2[1][2] = 2653ns;
slave_timing[3][160+19].t_rxd2[2][1] = 2750ns;

slave_timing[3][160+20].info_corner          = 2;
slave_timing[3][160+20].info_temp__j__       = -40;
slave_timing[3][160+20].info_i__quite_rec__  = 0.000000000;
slave_timing[3][160+20].info_dtr__ib__       = -1;
slave_timing[3][160+20].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+20].info_i__max_slave__  = 0.023000000;
slave_timing[3][160+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][160+20].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+20].t_rxd1[0][1] = 2814ns;
slave_timing[3][160+20].t_rxd1[1][0] = 2795ns;
slave_timing[3][160+20].t_rxd1[0][2] = 2115ns;
slave_timing[3][160+20].t_rxd1[2][0] = 3402ns;
slave_timing[3][160+20].t_rxd2[0][2] = 3330ns;
slave_timing[3][160+20].t_rxd2[2][0] = 2062ns;
slave_timing[3][160+20].t_rxd2[1][2] = 2779ns;
slave_timing[3][160+20].t_rxd2[2][1] = 2695ns;

slave_timing[3][160+21].info_corner          = 2;
slave_timing[3][160+21].info_temp__j__       = -40;
slave_timing[3][160+21].info_i__quite_rec__  = 0.000000000;
slave_timing[3][160+21].info_dtr__ib__       = -1;
slave_timing[3][160+21].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+21].info_i__max_slave__  = 0.025000000;
slave_timing[3][160+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][160+21].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+21].t_rxd1[0][1] = 2704ns;
slave_timing[3][160+21].t_rxd1[1][0] = 2880ns;
slave_timing[3][160+21].t_rxd1[0][2] = 2050ns;
slave_timing[3][160+21].t_rxd1[2][0] = 3457ns;
slave_timing[3][160+21].t_rxd2[0][2] = 3136ns;
slave_timing[3][160+21].t_rxd2[2][0] = 2204ns;
slave_timing[3][160+21].t_rxd2[1][2] = 2449ns;
slave_timing[3][160+21].t_rxd2[2][1] = 3024ns;

slave_timing[3][160+22].info_corner          = 2;
slave_timing[3][160+22].info_temp__j__       = -40;
slave_timing[3][160+22].info_i__quite_rec__  = 0.000000000;
slave_timing[3][160+22].info_dtr__ib__       = 1;
slave_timing[3][160+22].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+22].info_i__max_slave__  = 0.023000000;
slave_timing[3][160+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][160+22].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+22].t_rxd1[0][1] = 2896ns;
slave_timing[3][160+22].t_rxd1[1][0] = 2724ns;
slave_timing[3][160+22].t_rxd1[0][2] = 2156ns;
slave_timing[3][160+22].t_rxd1[2][0] = 3351ns;
slave_timing[3][160+22].t_rxd2[0][2] = 3501ns;
slave_timing[3][160+22].t_rxd2[2][0] = 1921ns;
slave_timing[3][160+22].t_rxd2[1][2] = 2989ns;
slave_timing[3][160+22].t_rxd2[2][1] = 2517ns;

slave_timing[3][160+23].info_corner          = 2;
slave_timing[3][160+23].info_temp__j__       = -40;
slave_timing[3][160+23].info_i__quite_rec__  = 0.000000000;
slave_timing[3][160+23].info_dtr__ib__       = 1;
slave_timing[3][160+23].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+23].info_i__max_slave__  = 0.025000000;
slave_timing[3][160+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][160+23].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+23].t_rxd1[0][1] = 2779ns;
slave_timing[3][160+23].t_rxd1[1][0] = 2811ns;
slave_timing[3][160+23].t_rxd1[0][2] = 2086ns;
slave_timing[3][160+23].t_rxd1[2][0] = 3407ns;
slave_timing[3][160+23].t_rxd2[0][2] = 3274ns;
slave_timing[3][160+23].t_rxd2[2][0] = 2095ns;
slave_timing[3][160+23].t_rxd2[1][2] = 2662ns;
slave_timing[3][160+23].t_rxd2[2][1] = 2755ns;

slave_timing[3][160+24].info_corner          = 2;
slave_timing[3][160+24].info_temp__j__       = -40;
slave_timing[3][160+24].info_i__quite_rec__  = 0.040000000;
slave_timing[3][160+24].info_dtr__ib__       = -1;
slave_timing[3][160+24].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+24].info_i__max_slave__  = 0.023000000;
slave_timing[3][160+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][160+24].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+24].t_rxd1[0][1] = 2742ns;
slave_timing[3][160+24].t_rxd1[1][0] = 2723ns;
slave_timing[3][160+24].t_rxd1[0][2] = 2024ns;
slave_timing[3][160+24].t_rxd1[2][0] = 3328ns;
slave_timing[3][160+24].t_rxd2[0][2] = 3288ns;
slave_timing[3][160+24].t_rxd2[2][0] = 2046ns;
slave_timing[3][160+24].t_rxd2[1][2] = 2732ns;
slave_timing[3][160+24].t_rxd2[2][1] = 2720ns;

slave_timing[3][160+25].info_corner          = 2;
slave_timing[3][160+25].info_temp__j__       = -40;
slave_timing[3][160+25].info_i__quite_rec__  = 0.040000000;
slave_timing[3][160+25].info_dtr__ib__       = -1;
slave_timing[3][160+25].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+25].info_i__max_slave__  = 0.025000000;
slave_timing[3][160+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][160+25].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+25].t_rxd1[0][1] = 2633ns;
slave_timing[3][160+25].t_rxd1[1][0] = 2808ns;
slave_timing[3][160+25].t_rxd1[0][2] = 1982ns;
slave_timing[3][160+25].t_rxd1[2][0] = 3379ns;
slave_timing[3][160+25].t_rxd2[0][2] = 3126ns;
slave_timing[3][160+25].t_rxd2[2][0] = 2190ns;
slave_timing[3][160+25].t_rxd2[1][2] = 2437ns;
slave_timing[3][160+25].t_rxd2[2][1] = 2970ns;

slave_timing[3][160+26].info_corner          = 2;
slave_timing[3][160+26].info_temp__j__       = -40;
slave_timing[3][160+26].info_i__quite_rec__  = 0.040000000;
slave_timing[3][160+26].info_dtr__ib__       = 1;
slave_timing[3][160+26].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+26].info_i__max_slave__  = 0.023000000;
slave_timing[3][160+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][160+26].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+26].t_rxd1[0][1] = 2807ns;
slave_timing[3][160+26].t_rxd1[1][0] = 2677ns;
slave_timing[3][160+26].t_rxd1[0][2] = 2086ns;
slave_timing[3][160+26].t_rxd1[2][0] = 3296ns;
slave_timing[3][160+26].t_rxd2[0][2] = 3479ns;
slave_timing[3][160+26].t_rxd2[2][0] = 1923ns;
slave_timing[3][160+26].t_rxd2[1][2] = 2963ns;
slave_timing[3][160+26].t_rxd2[2][1] = 2523ns;

slave_timing[3][160+27].info_corner          = 2;
slave_timing[3][160+27].info_temp__j__       = -40;
slave_timing[3][160+27].info_i__quite_rec__  = 0.040000000;
slave_timing[3][160+27].info_dtr__ib__       = 1;
slave_timing[3][160+27].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+27].info_i__max_slave__  = 0.025000000;
slave_timing[3][160+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][160+27].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+27].t_rxd1[0][1] = 2696ns;
slave_timing[3][160+27].t_rxd1[1][0] = 2762ns;
slave_timing[3][160+27].t_rxd1[0][2] = 2010ns;
slave_timing[3][160+27].t_rxd1[2][0] = 3350ns;
slave_timing[3][160+27].t_rxd2[0][2] = 3253ns;
slave_timing[3][160+27].t_rxd2[2][0] = 2090ns;
slave_timing[3][160+27].t_rxd2[1][2] = 2635ns;
slave_timing[3][160+27].t_rxd2[2][1] = 2809ns;

slave_timing[3][160+28].info_corner          = 2;
slave_timing[3][160+28].info_temp__j__       = -40;
slave_timing[3][160+28].info_i__quite_rec__  = 0.040000000;
slave_timing[3][160+28].info_dtr__ib__       = -1;
slave_timing[3][160+28].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+28].info_i__max_slave__  = 0.023000000;
slave_timing[3][160+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][160+28].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+28].t_rxd1[0][1] = 2775ns;
slave_timing[3][160+28].t_rxd1[1][0] = 2763ns;
slave_timing[3][160+28].t_rxd1[0][2] = 2081ns;
slave_timing[3][160+28].t_rxd1[2][0] = 3366ns;
slave_timing[3][160+28].t_rxd2[0][2] = 3330ns;
slave_timing[3][160+28].t_rxd2[2][0] = 2054ns;
slave_timing[3][160+28].t_rxd2[1][2] = 2737ns;
slave_timing[3][160+28].t_rxd2[2][1] = 2728ns;

slave_timing[3][160+29].info_corner          = 2;
slave_timing[3][160+29].info_temp__j__       = -40;
slave_timing[3][160+29].info_i__quite_rec__  = 0.040000000;
slave_timing[3][160+29].info_dtr__ib__       = -1;
slave_timing[3][160+29].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+29].info_i__max_slave__  = 0.025000000;
slave_timing[3][160+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][160+29].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+29].t_rxd1[0][1] = 2674ns;
slave_timing[3][160+29].t_rxd1[1][0] = 2842ns;
slave_timing[3][160+29].t_rxd1[0][2] = 2016ns;
slave_timing[3][160+29].t_rxd1[2][0] = 3419ns;
slave_timing[3][160+29].t_rxd2[0][2] = 3139ns;
slave_timing[3][160+29].t_rxd2[2][0] = 2196ns;
slave_timing[3][160+29].t_rxd2[1][2] = 2444ns;
slave_timing[3][160+29].t_rxd2[2][1] = 3015ns;

slave_timing[3][160+30].info_corner          = 2;
slave_timing[3][160+30].info_temp__j__       = -40;
slave_timing[3][160+30].info_i__quite_rec__  = 0.040000000;
slave_timing[3][160+30].info_dtr__ib__       = 1;
slave_timing[3][160+30].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+30].info_i__max_slave__  = 0.023000000;
slave_timing[3][160+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][160+30].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+30].t_rxd1[0][1] = 2845ns;
slave_timing[3][160+30].t_rxd1[1][0] = 2713ns;
slave_timing[3][160+30].t_rxd1[0][2] = 2113ns;
slave_timing[3][160+30].t_rxd1[2][0] = 3334ns;
slave_timing[3][160+30].t_rxd2[0][2] = 3489ns;
slave_timing[3][160+30].t_rxd2[2][0] = 1934ns;
slave_timing[3][160+30].t_rxd2[1][2] = 2974ns;
slave_timing[3][160+30].t_rxd2[2][1] = 2535ns;

slave_timing[3][160+31].info_corner          = 2;
slave_timing[3][160+31].info_temp__j__       = -40;
slave_timing[3][160+31].info_i__quite_rec__  = 0.040000000;
slave_timing[3][160+31].info_dtr__ib__       = 1;
slave_timing[3][160+31].info_i__offset_rec__ = 0.000000000;
slave_timing[3][160+31].info_i__max_slave__  = 0.025000000;
slave_timing[3][160+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][160+31].info_r__dsi_bus__    = 5.000;

slave_timing[3][160+31].t_rxd1[0][1] = 2731ns;
slave_timing[3][160+31].t_rxd1[1][0] = 2798ns;
slave_timing[3][160+31].t_rxd1[0][2] = 2053ns;
slave_timing[3][160+31].t_rxd1[2][0] = 3387ns;
slave_timing[3][160+31].t_rxd2[0][2] = 3265ns;
slave_timing[3][160+31].t_rxd2[2][0] = 2098ns;
slave_timing[3][160+31].t_rxd2[1][2] = 2645ns;
slave_timing[3][160+31].t_rxd2[2][1] = 2815ns;


slave_timing[1][128+0].info_corner          = 1;
slave_timing[1][128+0].info_temp__j__       = -40;
slave_timing[1][128+0].info_i__quite_rec__  = 0.006000000;
slave_timing[1][128+0].info_dtr__ib__       = -1;
slave_timing[1][128+0].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+0].info_i__max_slave__  = 0.023000000;
slave_timing[1][128+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][128+0].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+0].t_rxd1[0][1] = 1615ns;
slave_timing[1][128+0].t_rxd1[1][0] = 1639ns;
slave_timing[1][128+0].t_rxd1[0][2] = 1202ns;
slave_timing[1][128+0].t_rxd1[2][0] = 1986ns;
slave_timing[1][128+0].t_rxd2[0][2] = 1929ns;
slave_timing[1][128+0].t_rxd2[2][0] = 1229ns;
slave_timing[1][128+0].t_rxd2[1][2] = 1590ns;
slave_timing[1][128+0].t_rxd2[2][1] = 1631ns;

slave_timing[1][128+1].info_corner          = 1;
slave_timing[1][128+1].info_temp__j__       = -40;
slave_timing[1][128+1].info_i__quite_rec__  = 0.006000000;
slave_timing[1][128+1].info_dtr__ib__       = -1;
slave_timing[1][128+1].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+1].info_i__max_slave__  = 0.025000000;
slave_timing[1][128+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][128+1].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+1].t_rxd1[0][1] = 1556ns;
slave_timing[1][128+1].t_rxd1[1][0] = 1688ns;
slave_timing[1][128+1].t_rxd1[0][2] = 1185ns;
slave_timing[1][128+1].t_rxd1[2][0] = 2020ns;
slave_timing[1][128+1].t_rxd2[0][2] = 1834ns;
slave_timing[1][128+1].t_rxd2[2][0] = 1310ns;
slave_timing[1][128+1].t_rxd2[1][2] = 1423ns;
slave_timing[1][128+1].t_rxd2[2][1] = 1799ns;

slave_timing[1][128+2].info_corner          = 1;
slave_timing[1][128+2].info_temp__j__       = -40;
slave_timing[1][128+2].info_i__quite_rec__  = 0.006000000;
slave_timing[1][128+2].info_dtr__ib__       = 1;
slave_timing[1][128+2].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+2].info_i__max_slave__  = 0.023000000;
slave_timing[1][128+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][128+2].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+2].t_rxd1[0][1] = 1679ns;
slave_timing[1][128+2].t_rxd1[1][0] = 1593ns;
slave_timing[1][128+2].t_rxd1[0][2] = 1252ns;
slave_timing[1][128+2].t_rxd1[2][0] = 1953ns;
slave_timing[1][128+2].t_rxd2[0][2] = 2071ns;
slave_timing[1][128+2].t_rxd2[2][0] = 1145ns;
slave_timing[1][128+2].t_rxd2[1][2] = 1765ns;
slave_timing[1][128+2].t_rxd2[2][1] = 1484ns;

slave_timing[1][128+3].info_corner          = 1;
slave_timing[1][128+3].info_temp__j__       = -40;
slave_timing[1][128+3].info_i__quite_rec__  = 0.006000000;
slave_timing[1][128+3].info_dtr__ib__       = 1;
slave_timing[1][128+3].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+3].info_i__max_slave__  = 0.025000000;
slave_timing[1][128+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][128+3].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+3].t_rxd1[0][1] = 1611ns;
slave_timing[1][128+3].t_rxd1[1][0] = 1642ns;
slave_timing[1][128+3].t_rxd1[0][2] = 1216ns;
slave_timing[1][128+3].t_rxd1[2][0] = 1987ns;
slave_timing[1][128+3].t_rxd2[0][2] = 1930ns;
slave_timing[1][128+3].t_rxd2[2][0] = 1236ns;
slave_timing[1][128+3].t_rxd2[1][2] = 1570ns;
slave_timing[1][128+3].t_rxd2[2][1] = 1650ns;

slave_timing[1][128+4].info_corner          = 1;
slave_timing[1][128+4].info_temp__j__       = -40;
slave_timing[1][128+4].info_i__quite_rec__  = 0.006000000;
slave_timing[1][128+4].info_dtr__ib__       = -1;
slave_timing[1][128+4].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+4].info_i__max_slave__  = 0.023000000;
slave_timing[1][128+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][128+4].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+4].t_rxd1[0][1] = 1692ns;
slave_timing[1][128+4].t_rxd1[1][0] = 1711ns;
slave_timing[1][128+4].t_rxd1[0][2] = 1285ns;
slave_timing[1][128+4].t_rxd1[2][0] = 2055ns;
slave_timing[1][128+4].t_rxd2[0][2] = 1964ns;
slave_timing[1][128+4].t_rxd2[2][0] = 1247ns;
slave_timing[1][128+4].t_rxd2[1][2] = 1604ns;
slave_timing[1][128+4].t_rxd2[2][1] = 1644ns;

slave_timing[1][128+5].info_corner          = 1;
slave_timing[1][128+5].info_temp__j__       = -40;
slave_timing[1][128+5].info_i__quite_rec__  = 0.006000000;
slave_timing[1][128+5].info_dtr__ib__       = -1;
slave_timing[1][128+5].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+5].info_i__max_slave__  = 0.025000000;
slave_timing[1][128+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][128+5].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+5].t_rxd1[0][1] = 1628ns;
slave_timing[1][128+5].t_rxd1[1][0] = 1759ns;
slave_timing[1][128+5].t_rxd1[0][2] = 1249ns;
slave_timing[1][128+5].t_rxd1[2][0] = 2087ns;
slave_timing[1][128+5].t_rxd2[0][2] = 1852ns;
slave_timing[1][128+5].t_rxd2[2][0] = 1324ns;
slave_timing[1][128+5].t_rxd2[1][2] = 1437ns;
slave_timing[1][128+5].t_rxd2[2][1] = 1812ns;

slave_timing[1][128+6].info_corner          = 1;
slave_timing[1][128+6].info_temp__j__       = -40;
slave_timing[1][128+6].info_i__quite_rec__  = 0.006000000;
slave_timing[1][128+6].info_dtr__ib__       = 1;
slave_timing[1][128+6].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+6].info_i__max_slave__  = 0.023000000;
slave_timing[1][128+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][128+6].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+6].t_rxd1[0][1] = 1755ns;
slave_timing[1][128+6].t_rxd1[1][0] = 1662ns;
slave_timing[1][128+6].t_rxd1[0][2] = 1317ns;
slave_timing[1][128+6].t_rxd1[2][0] = 2022ns;
slave_timing[1][128+6].t_rxd2[0][2] = 2087ns;
slave_timing[1][128+6].t_rxd2[2][0] = 1162ns;
slave_timing[1][128+6].t_rxd2[1][2] = 1774ns;
slave_timing[1][128+6].t_rxd2[2][1] = 1497ns;

slave_timing[1][128+7].info_corner          = 1;
slave_timing[1][128+7].info_temp__j__       = -40;
slave_timing[1][128+7].info_i__quite_rec__  = 0.006000000;
slave_timing[1][128+7].info_dtr__ib__       = 1;
slave_timing[1][128+7].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+7].info_i__max_slave__  = 0.025000000;
slave_timing[1][128+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][128+7].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+7].t_rxd1[0][1] = 1684ns;
slave_timing[1][128+7].t_rxd1[1][0] = 1712ns;
slave_timing[1][128+7].t_rxd1[0][2] = 1279ns;
slave_timing[1][128+7].t_rxd1[2][0] = 2056ns;
slave_timing[1][128+7].t_rxd2[0][2] = 1947ns;
slave_timing[1][128+7].t_rxd2[2][0] = 1255ns;
slave_timing[1][128+7].t_rxd2[1][2] = 1584ns;
slave_timing[1][128+7].t_rxd2[2][1] = 1661ns;

slave_timing[1][128+8].info_corner          = 1;
slave_timing[1][128+8].info_temp__j__       = -40;
slave_timing[1][128+8].info_i__quite_rec__  = 0.003000000;
slave_timing[1][128+8].info_dtr__ib__       = -1;
slave_timing[1][128+8].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+8].info_i__max_slave__  = 0.023000000;
slave_timing[1][128+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][128+8].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+8].t_rxd1[0][1] = 1632ns;
slave_timing[1][128+8].t_rxd1[1][0] = 1626ns;
slave_timing[1][128+8].t_rxd1[0][2] = 1225ns;
slave_timing[1][128+8].t_rxd1[2][0] = 1975ns;
slave_timing[1][128+8].t_rxd2[0][2] = 1956ns;
slave_timing[1][128+8].t_rxd2[2][0] = 1220ns;
slave_timing[1][128+8].t_rxd2[1][2] = 1607ns;
slave_timing[1][128+8].t_rxd2[2][1] = 1620ns;

slave_timing[1][128+9].info_corner          = 1;
slave_timing[1][128+9].info_temp__j__       = -40;
slave_timing[1][128+9].info_i__quite_rec__  = 0.003000000;
slave_timing[1][128+9].info_dtr__ib__       = -1;
slave_timing[1][128+9].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+9].info_i__max_slave__  = 0.025000000;
slave_timing[1][128+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][128+9].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+9].t_rxd1[0][1] = 1569ns;
slave_timing[1][128+9].t_rxd1[1][0] = 1672ns;
slave_timing[1][128+9].t_rxd1[0][2] = 1193ns;
slave_timing[1][128+9].t_rxd1[2][0] = 2010ns;
slave_timing[1][128+9].t_rxd2[0][2] = 1842ns;
slave_timing[1][128+9].t_rxd2[2][0] = 1304ns;
slave_timing[1][128+9].t_rxd2[1][2] = 1438ns;
slave_timing[1][128+9].t_rxd2[2][1] = 1787ns;

slave_timing[1][128+10].info_corner          = 1;
slave_timing[1][128+10].info_temp__j__       = -40;
slave_timing[1][128+10].info_i__quite_rec__  = 0.003000000;
slave_timing[1][128+10].info_dtr__ib__       = 1;
slave_timing[1][128+10].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+10].info_i__max_slave__  = 0.023000000;
slave_timing[1][128+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][128+10].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+10].t_rxd1[0][1] = 1693ns;
slave_timing[1][128+10].t_rxd1[1][0] = 1573ns;
slave_timing[1][128+10].t_rxd1[0][2] = 1260ns;
slave_timing[1][128+10].t_rxd1[2][0] = 1939ns;
slave_timing[1][128+10].t_rxd2[0][2] = 2084ns;
slave_timing[1][128+10].t_rxd2[2][0] = 1140ns;
slave_timing[1][128+10].t_rxd2[1][2] = 1777ns;
slave_timing[1][128+10].t_rxd2[2][1] = 1470ns;

slave_timing[1][128+11].info_corner          = 1;
slave_timing[1][128+11].info_temp__j__       = -40;
slave_timing[1][128+11].info_i__quite_rec__  = 0.003000000;
slave_timing[1][128+11].info_dtr__ib__       = 1;
slave_timing[1][128+11].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+11].info_i__max_slave__  = 0.025000000;
slave_timing[1][128+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][128+11].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+11].t_rxd1[0][1] = 1624ns;
slave_timing[1][128+11].t_rxd1[1][0] = 1624ns;
slave_timing[1][128+11].t_rxd1[0][2] = 1221ns;
slave_timing[1][128+11].t_rxd1[2][0] = 1974ns;
slave_timing[1][128+11].t_rxd2[0][2] = 1938ns;
slave_timing[1][128+11].t_rxd2[2][0] = 1233ns;
slave_timing[1][128+11].t_rxd2[1][2] = 1586ns;
slave_timing[1][128+11].t_rxd2[2][1] = 1638ns;

slave_timing[1][128+12].info_corner          = 1;
slave_timing[1][128+12].info_temp__j__       = -40;
slave_timing[1][128+12].info_i__quite_rec__  = 0.003000000;
slave_timing[1][128+12].info_dtr__ib__       = -1;
slave_timing[1][128+12].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+12].info_i__max_slave__  = 0.023000000;
slave_timing[1][128+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][128+12].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+12].t_rxd1[0][1] = 1708ns;
slave_timing[1][128+12].t_rxd1[1][0] = 1696ns;
slave_timing[1][128+12].t_rxd1[0][2] = 1295ns;
slave_timing[1][128+12].t_rxd1[2][0] = 2045ns;
slave_timing[1][128+12].t_rxd2[0][2] = 1973ns;
slave_timing[1][128+12].t_rxd2[2][0] = 1240ns;
slave_timing[1][128+12].t_rxd2[1][2] = 1619ns;
slave_timing[1][128+12].t_rxd2[2][1] = 1630ns;

slave_timing[1][128+13].info_corner          = 1;
slave_timing[1][128+13].info_temp__j__       = -40;
slave_timing[1][128+13].info_i__quite_rec__  = 0.003000000;
slave_timing[1][128+13].info_dtr__ib__       = -1;
slave_timing[1][128+13].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+13].info_i__max_slave__  = 0.025000000;
slave_timing[1][128+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][128+13].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+13].t_rxd1[0][1] = 1645ns;
slave_timing[1][128+13].t_rxd1[1][0] = 1742ns;
slave_timing[1][128+13].t_rxd1[0][2] = 1259ns;
slave_timing[1][128+13].t_rxd1[2][0] = 2077ns;
slave_timing[1][128+13].t_rxd2[0][2] = 1860ns;
slave_timing[1][128+13].t_rxd2[2][0] = 1320ns;
slave_timing[1][128+13].t_rxd2[1][2] = 1451ns;
slave_timing[1][128+13].t_rxd2[2][1] = 1795ns;

slave_timing[1][128+14].info_corner          = 1;
slave_timing[1][128+14].info_temp__j__       = -40;
slave_timing[1][128+14].info_i__quite_rec__  = 0.003000000;
slave_timing[1][128+14].info_dtr__ib__       = 1;
slave_timing[1][128+14].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+14].info_i__max_slave__  = 0.023000000;
slave_timing[1][128+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][128+14].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+14].t_rxd1[0][1] = 1771ns;
slave_timing[1][128+14].t_rxd1[1][0] = 1646ns;
slave_timing[1][128+14].t_rxd1[0][2] = 1327ns;
slave_timing[1][128+14].t_rxd1[2][0] = 2007ns;
slave_timing[1][128+14].t_rxd2[0][2] = 2099ns;
slave_timing[1][128+14].t_rxd2[2][0] = 1156ns;
slave_timing[1][128+14].t_rxd2[1][2] = 1789ns;
slave_timing[1][128+14].t_rxd2[2][1] = 1484ns;

slave_timing[1][128+15].info_corner          = 1;
slave_timing[1][128+15].info_temp__j__       = -40;
slave_timing[1][128+15].info_i__quite_rec__  = 0.003000000;
slave_timing[1][128+15].info_dtr__ib__       = 1;
slave_timing[1][128+15].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+15].info_i__max_slave__  = 0.025000000;
slave_timing[1][128+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][128+15].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+15].t_rxd1[0][1] = 1701ns;
slave_timing[1][128+15].t_rxd1[1][0] = 1695ns;
slave_timing[1][128+15].t_rxd1[0][2] = 1290ns;
slave_timing[1][128+15].t_rxd1[2][0] = 2041ns;
slave_timing[1][128+15].t_rxd2[0][2] = 1956ns;
slave_timing[1][128+15].t_rxd2[2][0] = 1248ns;
slave_timing[1][128+15].t_rxd2[1][2] = 1595ns;
slave_timing[1][128+15].t_rxd2[2][1] = 1646ns;

slave_timing[1][128+16].info_corner          = 1;
slave_timing[1][128+16].info_temp__j__       = -40;
slave_timing[1][128+16].info_i__quite_rec__  = 0.000000000;
slave_timing[1][128+16].info_dtr__ib__       = -1;
slave_timing[1][128+16].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+16].info_i__max_slave__  = 0.023000000;
slave_timing[1][128+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][128+16].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+16].t_rxd1[0][1] = 1622ns;
slave_timing[1][128+16].t_rxd1[1][0] = 1629ns;
slave_timing[1][128+16].t_rxd1[0][2] = 1219ns;
slave_timing[1][128+16].t_rxd1[2][0] = 1981ns;
slave_timing[1][128+16].t_rxd2[0][2] = 1950ns;
slave_timing[1][128+16].t_rxd2[2][0] = 1228ns;
slave_timing[1][128+16].t_rxd2[1][2] = 1599ns;
slave_timing[1][128+16].t_rxd2[2][1] = 1629ns;

slave_timing[1][128+17].info_corner          = 1;
slave_timing[1][128+17].info_temp__j__       = -40;
slave_timing[1][128+17].info_i__quite_rec__  = 0.000000000;
slave_timing[1][128+17].info_dtr__ib__       = -1;
slave_timing[1][128+17].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+17].info_i__max_slave__  = 0.025000000;
slave_timing[1][128+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][128+17].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+17].t_rxd1[0][1] = 1561ns;
slave_timing[1][128+17].t_rxd1[1][0] = 1681ns;
slave_timing[1][128+17].t_rxd1[0][2] = 1188ns;
slave_timing[1][128+17].t_rxd1[2][0] = 2015ns;
slave_timing[1][128+17].t_rxd2[0][2] = 1836ns;
slave_timing[1][128+17].t_rxd2[2][0] = 1308ns;
slave_timing[1][128+17].t_rxd2[1][2] = 1427ns;
slave_timing[1][128+17].t_rxd2[2][1] = 1800ns;

slave_timing[1][128+18].info_corner          = 1;
slave_timing[1][128+18].info_temp__j__       = -40;
slave_timing[1][128+18].info_i__quite_rec__  = 0.000000000;
slave_timing[1][128+18].info_dtr__ib__       = 1;
slave_timing[1][128+18].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+18].info_i__max_slave__  = 0.023000000;
slave_timing[1][128+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][128+18].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+18].t_rxd1[0][1] = 1682ns;
slave_timing[1][128+18].t_rxd1[1][0] = 1589ns;
slave_timing[1][128+18].t_rxd1[0][2] = 1252ns;
slave_timing[1][128+18].t_rxd1[2][0] = 1949ns;
slave_timing[1][128+18].t_rxd2[0][2] = 2071ns;
slave_timing[1][128+18].t_rxd2[2][0] = 1141ns;
slave_timing[1][128+18].t_rxd2[1][2] = 1768ns;
slave_timing[1][128+18].t_rxd2[2][1] = 1474ns;

slave_timing[1][128+19].info_corner          = 1;
slave_timing[1][128+19].info_temp__j__       = -40;
slave_timing[1][128+19].info_i__quite_rec__  = 0.000000000;
slave_timing[1][128+19].info_dtr__ib__       = 1;
slave_timing[1][128+19].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+19].info_i__max_slave__  = 0.025000000;
slave_timing[1][128+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][128+19].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+19].t_rxd1[0][1] = 1612ns;
slave_timing[1][128+19].t_rxd1[1][0] = 1638ns;
slave_timing[1][128+19].t_rxd1[0][2] = 1214ns;
slave_timing[1][128+19].t_rxd1[2][0] = 1985ns;
slave_timing[1][128+19].t_rxd2[0][2] = 1929ns;
slave_timing[1][128+19].t_rxd2[2][0] = 1234ns;
slave_timing[1][128+19].t_rxd2[1][2] = 1571ns;
slave_timing[1][128+19].t_rxd2[2][1] = 1644ns;

slave_timing[1][128+20].info_corner          = 1;
slave_timing[1][128+20].info_temp__j__       = -40;
slave_timing[1][128+20].info_i__quite_rec__  = 0.000000000;
slave_timing[1][128+20].info_dtr__ib__       = -1;
slave_timing[1][128+20].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+20].info_i__max_slave__  = 0.023000000;
slave_timing[1][128+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][128+20].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+20].t_rxd1[0][1] = 1700ns;
slave_timing[1][128+20].t_rxd1[1][0] = 1702ns;
slave_timing[1][128+20].t_rxd1[0][2] = 1288ns;
slave_timing[1][128+20].t_rxd1[2][0] = 2048ns;
slave_timing[1][128+20].t_rxd2[0][2] = 1966ns;
slave_timing[1][128+20].t_rxd2[2][0] = 1244ns;
slave_timing[1][128+20].t_rxd2[1][2] = 1607ns;
slave_timing[1][128+20].t_rxd2[2][1] = 1638ns;

slave_timing[1][128+21].info_corner          = 1;
slave_timing[1][128+21].info_temp__j__       = -40;
slave_timing[1][128+21].info_i__quite_rec__  = 0.000000000;
slave_timing[1][128+21].info_dtr__ib__       = -1;
slave_timing[1][128+21].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+21].info_i__max_slave__  = 0.025000000;
slave_timing[1][128+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][128+21].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+21].t_rxd1[0][1] = 1635ns;
slave_timing[1][128+21].t_rxd1[1][0] = 1750ns;
slave_timing[1][128+21].t_rxd1[0][2] = 1254ns;
slave_timing[1][128+21].t_rxd1[2][0] = 2082ns;
slave_timing[1][128+21].t_rxd2[0][2] = 1854ns;
slave_timing[1][128+21].t_rxd2[2][0] = 1324ns;
slave_timing[1][128+21].t_rxd2[1][2] = 1438ns;
slave_timing[1][128+21].t_rxd2[2][1] = 1808ns;

slave_timing[1][128+22].info_corner          = 1;
slave_timing[1][128+22].info_temp__j__       = -40;
slave_timing[1][128+22].info_i__quite_rec__  = 0.000000000;
slave_timing[1][128+22].info_dtr__ib__       = 1;
slave_timing[1][128+22].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+22].info_i__max_slave__  = 0.023000000;
slave_timing[1][128+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][128+22].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+22].t_rxd1[0][1] = 1760ns;
slave_timing[1][128+22].t_rxd1[1][0] = 1657ns;
slave_timing[1][128+22].t_rxd1[0][2] = 1319ns;
slave_timing[1][128+22].t_rxd1[2][0] = 2018ns;
slave_timing[1][128+22].t_rxd2[0][2] = 2086ns;
slave_timing[1][128+22].t_rxd2[2][0] = 1160ns;
slave_timing[1][128+22].t_rxd2[1][2] = 1777ns;
slave_timing[1][128+22].t_rxd2[2][1] = 1491ns;

slave_timing[1][128+23].info_corner          = 1;
slave_timing[1][128+23].info_temp__j__       = -40;
slave_timing[1][128+23].info_i__quite_rec__  = 0.000000000;
slave_timing[1][128+23].info_dtr__ib__       = 1;
slave_timing[1][128+23].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+23].info_i__max_slave__  = 0.025000000;
slave_timing[1][128+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][128+23].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+23].t_rxd1[0][1] = 1688ns;
slave_timing[1][128+23].t_rxd1[1][0] = 1708ns;
slave_timing[1][128+23].t_rxd1[0][2] = 1283ns;
slave_timing[1][128+23].t_rxd1[2][0] = 2051ns;
slave_timing[1][128+23].t_rxd2[0][2] = 1947ns;
slave_timing[1][128+23].t_rxd2[2][0] = 1250ns;
slave_timing[1][128+23].t_rxd2[1][2] = 1583ns;
slave_timing[1][128+23].t_rxd2[2][1] = 1656ns;

slave_timing[1][128+24].info_corner          = 1;
slave_timing[1][128+24].info_temp__j__       = -40;
slave_timing[1][128+24].info_i__quite_rec__  = 0.040000000;
slave_timing[1][128+24].info_dtr__ib__       = -1;
slave_timing[1][128+24].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+24].info_i__max_slave__  = 0.023000000;
slave_timing[1][128+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][128+24].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+24].t_rxd1[0][1] = 1624ns;
slave_timing[1][128+24].t_rxd1[1][0] = 1610ns;
slave_timing[1][128+24].t_rxd1[0][2] = 1223ns;
slave_timing[1][128+24].t_rxd1[2][0] = 1962ns;
slave_timing[1][128+24].t_rxd2[0][2] = 1957ns;
slave_timing[1][128+24].t_rxd2[2][0] = 1219ns;
slave_timing[1][128+24].t_rxd2[1][2] = 1611ns;
slave_timing[1][128+24].t_rxd2[2][1] = 1616ns;

slave_timing[1][128+25].info_corner          = 1;
slave_timing[1][128+25].info_temp__j__       = -40;
slave_timing[1][128+25].info_i__quite_rec__  = 0.040000000;
slave_timing[1][128+25].info_dtr__ib__       = -1;
slave_timing[1][128+25].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+25].info_i__max_slave__  = 0.025000000;
slave_timing[1][128+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][128+25].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+25].t_rxd1[0][1] = 1565ns;
slave_timing[1][128+25].t_rxd1[1][0] = 1659ns;
slave_timing[1][128+25].t_rxd1[0][2] = 1185ns;
slave_timing[1][128+25].t_rxd1[2][0] = 1995ns;
slave_timing[1][128+25].t_rxd2[0][2] = 1842ns;
slave_timing[1][128+25].t_rxd2[2][0] = 1300ns;
slave_timing[1][128+25].t_rxd2[1][2] = 1443ns;
slave_timing[1][128+25].t_rxd2[2][1] = 1784ns;

slave_timing[1][128+26].info_corner          = 1;
slave_timing[1][128+26].info_temp__j__       = -40;
slave_timing[1][128+26].info_i__quite_rec__  = 0.040000000;
slave_timing[1][128+26].info_dtr__ib__       = 1;
slave_timing[1][128+26].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+26].info_i__max_slave__  = 0.023000000;
slave_timing[1][128+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][128+26].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+26].t_rxd1[0][1] = 1669ns;
slave_timing[1][128+26].t_rxd1[1][0] = 1584ns;
slave_timing[1][128+26].t_rxd1[0][2] = 1242ns;
slave_timing[1][128+26].t_rxd1[2][0] = 1943ns;
slave_timing[1][128+26].t_rxd2[0][2] = 2069ns;
slave_timing[1][128+26].t_rxd2[2][0] = 1148ns;
slave_timing[1][128+26].t_rxd2[1][2] = 1762ns;
slave_timing[1][128+26].t_rxd2[2][1] = 1488ns;

slave_timing[1][128+27].info_corner          = 1;
slave_timing[1][128+27].info_temp__j__       = -40;
slave_timing[1][128+27].info_i__quite_rec__  = 0.040000000;
slave_timing[1][128+27].info_dtr__ib__       = 1;
slave_timing[1][128+27].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+27].info_i__max_slave__  = 0.025000000;
slave_timing[1][128+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][128+27].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+27].t_rxd1[0][1] = 1600ns;
slave_timing[1][128+27].t_rxd1[1][0] = 1632ns;
slave_timing[1][128+27].t_rxd1[0][2] = 1207ns;
slave_timing[1][128+27].t_rxd1[2][0] = 1976ns;
slave_timing[1][128+27].t_rxd2[0][2] = 1929ns;
slave_timing[1][128+27].t_rxd2[2][0] = 1241ns;
slave_timing[1][128+27].t_rxd2[1][2] = 1566ns;
slave_timing[1][128+27].t_rxd2[2][1] = 1656ns;

slave_timing[1][128+28].info_corner          = 1;
slave_timing[1][128+28].info_temp__j__       = -40;
slave_timing[1][128+28].info_i__quite_rec__  = 0.040000000;
slave_timing[1][128+28].info_dtr__ib__       = -1;
slave_timing[1][128+28].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+28].info_i__max_slave__  = 0.023000000;
slave_timing[1][128+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][128+28].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+28].t_rxd1[0][1] = 1668ns;
slave_timing[1][128+28].t_rxd1[1][0] = 1650ns;
slave_timing[1][128+28].t_rxd1[0][2] = 1261ns;
slave_timing[1][128+28].t_rxd1[2][0] = 2002ns;
slave_timing[1][128+28].t_rxd2[0][2] = 1970ns;
slave_timing[1][128+28].t_rxd2[2][0] = 1236ns;
slave_timing[1][128+28].t_rxd2[1][2] = 1622ns;
slave_timing[1][128+28].t_rxd2[2][1] = 1629ns;

slave_timing[1][128+29].info_corner          = 1;
slave_timing[1][128+29].info_temp__j__       = -40;
slave_timing[1][128+29].info_i__quite_rec__  = 0.040000000;
slave_timing[1][128+29].info_dtr__ib__       = -1;
slave_timing[1][128+29].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+29].info_i__max_slave__  = 0.025000000;
slave_timing[1][128+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][128+29].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+29].t_rxd1[0][1] = 1604ns;
slave_timing[1][128+29].t_rxd1[1][0] = 1703ns;
slave_timing[1][128+29].t_rxd1[0][2] = 1225ns;
slave_timing[1][128+29].t_rxd1[2][0] = 2037ns;
slave_timing[1][128+29].t_rxd2[0][2] = 1855ns;
slave_timing[1][128+29].t_rxd2[2][0] = 1318ns;
slave_timing[1][128+29].t_rxd2[1][2] = 1453ns;
slave_timing[1][128+29].t_rxd2[2][1] = 1795ns;

slave_timing[1][128+30].info_corner          = 1;
slave_timing[1][128+30].info_temp__j__       = -40;
slave_timing[1][128+30].info_i__quite_rec__  = 0.040000000;
slave_timing[1][128+30].info_dtr__ib__       = 1;
slave_timing[1][128+30].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+30].info_i__max_slave__  = 0.023000000;
slave_timing[1][128+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][128+30].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+30].t_rxd1[0][1] = 1710ns;
slave_timing[1][128+30].t_rxd1[1][0] = 1627ns;
slave_timing[1][128+30].t_rxd1[0][2] = 1282ns;
slave_timing[1][128+30].t_rxd1[2][0] = 1986ns;
slave_timing[1][128+30].t_rxd2[0][2] = 2081ns;
slave_timing[1][128+30].t_rxd2[2][0] = 1165ns;
slave_timing[1][128+30].t_rxd2[1][2] = 1771ns;
slave_timing[1][128+30].t_rxd2[2][1] = 1502ns;

slave_timing[1][128+31].info_corner          = 1;
slave_timing[1][128+31].info_temp__j__       = -40;
slave_timing[1][128+31].info_i__quite_rec__  = 0.040000000;
slave_timing[1][128+31].info_dtr__ib__       = 1;
slave_timing[1][128+31].info_i__offset_rec__ = 0.000000000;
slave_timing[1][128+31].info_i__max_slave__  = 0.025000000;
slave_timing[1][128+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][128+31].info_r__dsi_bus__    = 5.000;

slave_timing[1][128+31].t_rxd1[0][1] = 1642ns;
slave_timing[1][128+31].t_rxd1[1][0] = 1674ns;
slave_timing[1][128+31].t_rxd1[0][2] = 1246ns;
slave_timing[1][128+31].t_rxd1[2][0] = 2019ns;
slave_timing[1][128+31].t_rxd2[0][2] = 1940ns;
slave_timing[1][128+31].t_rxd2[2][0] = 1256ns;
slave_timing[1][128+31].t_rxd2[1][2] = 1576ns;
slave_timing[1][128+31].t_rxd2[2][1] = 1663ns;

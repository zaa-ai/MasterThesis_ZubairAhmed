/* ###   interface instances   ###################################################### */

SRAM_BIST_registers_SRAM_ECC_CONTROL_if SRAM_BIST_registers_SRAM_ECC_CONTROL (); 
SRAM_BIST_registers_SRAM_BIST_CTRL_if SRAM_BIST_registers_SRAM_BIST_CTRL (); 
SRAM_BIST_registers_SRAM_BIST_STAT_if SRAM_BIST_registers_SRAM_BIST_STAT (); 



slave_timing[3][32+0].info_corner          = 2;
slave_timing[3][32+0].info_temp__j__       = 125;
slave_timing[3][32+0].info_i__quite_rec__  = 0.006000000;
slave_timing[3][32+0].info_dtr__ib__       = -1;
slave_timing[3][32+0].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+0].info_i__max_slave__  = 0.023000000;
slave_timing[3][32+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][32+0].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+0].t_rxd1[0][1] = 2760ns;
slave_timing[3][32+0].t_rxd1[1][0] = 2767ns;
slave_timing[3][32+0].t_rxd1[0][2] = 2068ns;
slave_timing[3][32+0].t_rxd1[2][0] = 3355ns;
slave_timing[3][32+0].t_rxd2[0][2] = 3326ns;
slave_timing[3][32+0].t_rxd2[2][0] = 2065ns;
slave_timing[3][32+0].t_rxd2[1][2] = 2750ns;
slave_timing[3][32+0].t_rxd2[2][1] = 2747ns;

slave_timing[3][32+1].info_corner          = 2;
slave_timing[3][32+1].info_temp__j__       = 125;
slave_timing[3][32+1].info_i__quite_rec__  = 0.006000000;
slave_timing[3][32+1].info_dtr__ib__       = -1;
slave_timing[3][32+1].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+1].info_i__max_slave__  = 0.025000000;
slave_timing[3][32+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][32+1].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+1].t_rxd1[0][1] = 2656ns;
slave_timing[3][32+1].t_rxd1[1][0] = 2850ns;
slave_timing[3][32+1].t_rxd1[0][2] = 2007ns;
slave_timing[3][32+1].t_rxd1[2][0] = 3409ns;
slave_timing[3][32+1].t_rxd2[0][2] = 3138ns;
slave_timing[3][32+1].t_rxd2[2][0] = 2219ns;
slave_timing[3][32+1].t_rxd2[1][2] = 2465ns;
slave_timing[3][32+1].t_rxd2[2][1] = 3031ns;

slave_timing[3][32+2].info_corner          = 2;
slave_timing[3][32+2].info_temp__j__       = 125;
slave_timing[3][32+2].info_i__quite_rec__  = 0.006000000;
slave_timing[3][32+2].info_dtr__ib__       = 1;
slave_timing[3][32+2].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+2].info_i__max_slave__  = 0.023000000;
slave_timing[3][32+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][32+2].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+2].t_rxd1[0][1] = 2825ns;
slave_timing[3][32+2].t_rxd1[1][0] = 2703ns;
slave_timing[3][32+2].t_rxd1[0][2] = 2094ns;
slave_timing[3][32+2].t_rxd1[2][0] = 3304ns;
slave_timing[3][32+2].t_rxd2[0][2] = 3493ns;
slave_timing[3][32+2].t_rxd2[2][0] = 1929ns;
slave_timing[3][32+2].t_rxd2[1][2] = 3003ns;
slave_timing[3][32+2].t_rxd2[2][1] = 2521ns;

slave_timing[3][32+3].info_corner          = 2;
slave_timing[3][32+3].info_temp__j__       = 125;
slave_timing[3][32+3].info_i__quite_rec__  = 0.006000000;
slave_timing[3][32+3].info_dtr__ib__       = 1;
slave_timing[3][32+3].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+3].info_i__max_slave__  = 0.025000000;
slave_timing[3][32+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][32+3].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+3].t_rxd1[0][1] = 2709ns;
slave_timing[3][32+3].t_rxd1[1][0] = 2783ns;
slave_timing[3][32+3].t_rxd1[0][2] = 2025ns;
slave_timing[3][32+3].t_rxd1[2][0] = 3357ns;
slave_timing[3][32+3].t_rxd2[0][2] = 3266ns;
slave_timing[3][32+3].t_rxd2[2][0] = 2098ns;
slave_timing[3][32+3].t_rxd2[1][2] = 2670ns;
slave_timing[3][32+3].t_rxd2[2][1] = 2804ns;

slave_timing[3][32+4].info_corner          = 2;
slave_timing[3][32+4].info_temp__j__       = 125;
slave_timing[3][32+4].info_i__quite_rec__  = 0.006000000;
slave_timing[3][32+4].info_dtr__ib__       = -1;
slave_timing[3][32+4].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+4].info_i__max_slave__  = 0.023000000;
slave_timing[3][32+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][32+4].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+4].t_rxd1[0][1] = 2913ns;
slave_timing[3][32+4].t_rxd1[1][0] = 2908ns;
slave_timing[3][32+4].t_rxd1[0][2] = 2210ns;
slave_timing[3][32+4].t_rxd1[2][0] = 3488ns;
slave_timing[3][32+4].t_rxd2[0][2] = 3348ns;
slave_timing[3][32+4].t_rxd2[2][0] = 2094ns;
slave_timing[3][32+4].t_rxd2[1][2] = 2771ns;
slave_timing[3][32+4].t_rxd2[2][1] = 2766ns;

slave_timing[3][32+5].info_corner          = 2;
slave_timing[3][32+5].info_temp__j__       = 125;
slave_timing[3][32+5].info_i__quite_rec__  = 0.006000000;
slave_timing[3][32+5].info_dtr__ib__       = -1;
slave_timing[3][32+5].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+5].info_i__max_slave__  = 0.025000000;
slave_timing[3][32+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][32+5].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+5].t_rxd1[0][1] = 2806ns;
slave_timing[3][32+5].t_rxd1[1][0] = 2989ns;
slave_timing[3][32+5].t_rxd1[0][2] = 2146ns;
slave_timing[3][32+5].t_rxd1[2][0] = 3540ns;
slave_timing[3][32+5].t_rxd2[0][2] = 3160ns;
slave_timing[3][32+5].t_rxd2[2][0] = 2242ns;
slave_timing[3][32+5].t_rxd2[1][2] = 2487ns;
slave_timing[3][32+5].t_rxd2[2][1] = 3052ns;

slave_timing[3][32+6].info_corner          = 2;
slave_timing[3][32+6].info_temp__j__       = 125;
slave_timing[3][32+6].info_i__quite_rec__  = 0.006000000;
slave_timing[3][32+6].info_dtr__ib__       = 1;
slave_timing[3][32+6].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+6].info_i__max_slave__  = 0.023000000;
slave_timing[3][32+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][32+6].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+6].t_rxd1[0][1] = 2985ns;
slave_timing[3][32+6].t_rxd1[1][0] = 2835ns;
slave_timing[3][32+6].t_rxd1[0][2] = 2239ns;
slave_timing[3][32+6].t_rxd1[2][0] = 3433ns;
slave_timing[3][32+6].t_rxd2[0][2] = 3516ns;
slave_timing[3][32+6].t_rxd2[2][0] = 1950ns;
slave_timing[3][32+6].t_rxd2[1][2] = 3070ns;
slave_timing[3][32+6].t_rxd2[2][1] = 2503ns;

slave_timing[3][32+7].info_corner          = 2;
slave_timing[3][32+7].info_temp__j__       = 125;
slave_timing[3][32+7].info_i__quite_rec__  = 0.006000000;
slave_timing[3][32+7].info_dtr__ib__       = 1;
slave_timing[3][32+7].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+7].info_i__max_slave__  = 0.025000000;
slave_timing[3][32+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][32+7].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+7].t_rxd1[0][1] = 2912ns;
slave_timing[3][32+7].t_rxd1[1][0] = 2922ns;
slave_timing[3][32+7].t_rxd1[0][2] = 2175ns;
slave_timing[3][32+7].t_rxd1[2][0] = 3488ns;
slave_timing[3][32+7].t_rxd2[0][2] = 3288ns;
slave_timing[3][32+7].t_rxd2[2][0] = 2119ns;
slave_timing[3][32+7].t_rxd2[1][2] = 2728ns;
slave_timing[3][32+7].t_rxd2[2][1] = 2785ns;

slave_timing[3][32+8].info_corner          = 2;
slave_timing[3][32+8].info_temp__j__       = 125;
slave_timing[3][32+8].info_i__quite_rec__  = 0.003000000;
slave_timing[3][32+8].info_dtr__ib__       = -1;
slave_timing[3][32+8].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+8].info_i__max_slave__  = 0.023000000;
slave_timing[3][32+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][32+8].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+8].t_rxd1[0][1] = 2752ns;
slave_timing[3][32+8].t_rxd1[1][0] = 2740ns;
slave_timing[3][32+8].t_rxd1[0][2] = 2054ns;
slave_timing[3][32+8].t_rxd1[2][0] = 3326ns;
slave_timing[3][32+8].t_rxd2[0][2] = 3325ns;
slave_timing[3][32+8].t_rxd2[2][0] = 2041ns;
slave_timing[3][32+8].t_rxd2[1][2] = 2766ns;
slave_timing[3][32+8].t_rxd2[2][1] = 2674ns;

slave_timing[3][32+9].info_corner          = 2;
slave_timing[3][32+9].info_temp__j__       = 125;
slave_timing[3][32+9].info_i__quite_rec__  = 0.003000000;
slave_timing[3][32+9].info_dtr__ib__       = -1;
slave_timing[3][32+9].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+9].info_i__max_slave__  = 0.025000000;
slave_timing[3][32+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][32+9].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+9].t_rxd1[0][1] = 2648ns;
slave_timing[3][32+9].t_rxd1[1][0] = 2820ns;
slave_timing[3][32+9].t_rxd1[0][2] = 1987ns;
slave_timing[3][32+9].t_rxd1[2][0] = 3381ns;
slave_timing[3][32+9].t_rxd2[0][2] = 3129ns;
slave_timing[3][32+9].t_rxd2[2][0] = 2192ns;
slave_timing[3][32+9].t_rxd2[1][2] = 2473ns;
slave_timing[3][32+9].t_rxd2[2][1] = 2987ns;

slave_timing[3][32+10].info_corner          = 2;
slave_timing[3][32+10].info_temp__j__       = 125;
slave_timing[3][32+10].info_i__quite_rec__  = 0.003000000;
slave_timing[3][32+10].info_dtr__ib__       = 1;
slave_timing[3][32+10].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+10].info_i__max_slave__  = 0.023000000;
slave_timing[3][32+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][32+10].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+10].t_rxd1[0][1] = 2814ns;
slave_timing[3][32+10].t_rxd1[1][0] = 2644ns;
slave_timing[3][32+10].t_rxd1[0][2] = 2080ns;
slave_timing[3][32+10].t_rxd1[2][0] = 3255ns;
slave_timing[3][32+10].t_rxd2[0][2] = 3493ns;
slave_timing[3][32+10].t_rxd2[2][0] = 1906ns;
slave_timing[3][32+10].t_rxd2[1][2] = 3006ns;
slave_timing[3][32+10].t_rxd2[2][1] = 2492ns;

slave_timing[3][32+11].info_corner          = 2;
slave_timing[3][32+11].info_temp__j__       = 125;
slave_timing[3][32+11].info_i__quite_rec__  = 0.003000000;
slave_timing[3][32+11].info_dtr__ib__       = 1;
slave_timing[3][32+11].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+11].info_i__max_slave__  = 0.025000000;
slave_timing[3][32+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][32+11].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+11].t_rxd1[0][1] = 2695ns;
slave_timing[3][32+11].t_rxd1[1][0] = 2725ns;
slave_timing[3][32+11].t_rxd1[0][2] = 2015ns;
slave_timing[3][32+11].t_rxd1[2][0] = 3308ns;
slave_timing[3][32+11].t_rxd2[0][2] = 3260ns;
slave_timing[3][32+11].t_rxd2[2][0] = 2082ns;
slave_timing[3][32+11].t_rxd2[1][2] = 2671ns;
slave_timing[3][32+11].t_rxd2[2][1] = 2774ns;

slave_timing[3][32+12].info_corner          = 2;
slave_timing[3][32+12].info_temp__j__       = 125;
slave_timing[3][32+12].info_i__quite_rec__  = 0.003000000;
slave_timing[3][32+12].info_dtr__ib__       = -1;
slave_timing[3][32+12].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+12].info_i__max_slave__  = 0.023000000;
slave_timing[3][32+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][32+12].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+12].t_rxd1[0][1] = 2925ns;
slave_timing[3][32+12].t_rxd1[1][0] = 2879ns;
slave_timing[3][32+12].t_rxd1[0][2] = 2212ns;
slave_timing[3][32+12].t_rxd1[2][0] = 3455ns;
slave_timing[3][32+12].t_rxd2[0][2] = 3348ns;
slave_timing[3][32+12].t_rxd2[2][0] = 2073ns;
slave_timing[3][32+12].t_rxd2[1][2] = 2787ns;
slave_timing[3][32+12].t_rxd2[2][1] = 2732ns;

slave_timing[3][32+13].info_corner          = 2;
slave_timing[3][32+13].info_temp__j__       = 125;
slave_timing[3][32+13].info_i__quite_rec__  = 0.003000000;
slave_timing[3][32+13].info_dtr__ib__       = -1;
slave_timing[3][32+13].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+13].info_i__max_slave__  = 0.025000000;
slave_timing[3][32+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][32+13].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+13].t_rxd1[0][1] = 2811ns;
slave_timing[3][32+13].t_rxd1[1][0] = 2961ns;
slave_timing[3][32+13].t_rxd1[0][2] = 2143ns;
slave_timing[3][32+13].t_rxd1[2][0] = 3510ns;
slave_timing[3][32+13].t_rxd2[0][2] = 3154ns;
slave_timing[3][32+13].t_rxd2[2][0] = 2222ns;
slave_timing[3][32+13].t_rxd2[1][2] = 2499ns;
slave_timing[3][32+13].t_rxd2[2][1] = 3010ns;

slave_timing[3][32+14].info_corner          = 2;
slave_timing[3][32+14].info_temp__j__       = 125;
slave_timing[3][32+14].info_i__quite_rec__  = 0.003000000;
slave_timing[3][32+14].info_dtr__ib__       = 1;
slave_timing[3][32+14].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+14].info_i__max_slave__  = 0.023000000;
slave_timing[3][32+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][32+14].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+14].t_rxd1[0][1] = 2981ns;
slave_timing[3][32+14].t_rxd1[1][0] = 2790ns;
slave_timing[3][32+14].t_rxd1[0][2] = 2238ns;
slave_timing[3][32+14].t_rxd1[2][0] = 3380ns;
slave_timing[3][32+14].t_rxd2[0][2] = 3508ns;
slave_timing[3][32+14].t_rxd2[2][0] = 1931ns;
slave_timing[3][32+14].t_rxd2[1][2] = 3026ns;
slave_timing[3][32+14].t_rxd2[2][1] = 2517ns;

slave_timing[3][32+15].info_corner          = 2;
slave_timing[3][32+15].info_temp__j__       = 125;
slave_timing[3][32+15].info_i__quite_rec__  = 0.003000000;
slave_timing[3][32+15].info_dtr__ib__       = 1;
slave_timing[3][32+15].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+15].info_i__max_slave__  = 0.025000000;
slave_timing[3][32+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][32+15].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+15].t_rxd1[0][1] = 2862ns;
slave_timing[3][32+15].t_rxd1[1][0] = 2868ns;
slave_timing[3][32+15].t_rxd1[0][2] = 2171ns;
slave_timing[3][32+15].t_rxd1[2][0] = 3436ns;
slave_timing[3][32+15].t_rxd2[0][2] = 3278ns;
slave_timing[3][32+15].t_rxd2[2][0] = 2101ns;
slave_timing[3][32+15].t_rxd2[1][2] = 2694ns;
slave_timing[3][32+15].t_rxd2[2][1] = 2793ns;

slave_timing[3][32+16].info_corner          = 2;
slave_timing[3][32+16].info_temp__j__       = 125;
slave_timing[3][32+16].info_i__quite_rec__  = 0.000000000;
slave_timing[3][32+16].info_dtr__ib__       = -1;
slave_timing[3][32+16].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+16].info_i__max_slave__  = 0.023000000;
slave_timing[3][32+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][32+16].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+16].t_rxd1[0][1] = 2731ns;
slave_timing[3][32+16].t_rxd1[1][0] = 2689ns;
slave_timing[3][32+16].t_rxd1[0][2] = 2037ns;
slave_timing[3][32+16].t_rxd1[2][0] = 3280ns;
slave_timing[3][32+16].t_rxd2[0][2] = 3313ns;
slave_timing[3][32+16].t_rxd2[2][0] = 2025ns;
slave_timing[3][32+16].t_rxd2[1][2] = 2761ns;
slave_timing[3][32+16].t_rxd2[2][1] = 2687ns;

slave_timing[3][32+17].info_corner          = 2;
slave_timing[3][32+17].info_temp__j__       = 125;
slave_timing[3][32+17].info_i__quite_rec__  = 0.000000000;
slave_timing[3][32+17].info_dtr__ib__       = -1;
slave_timing[3][32+17].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+17].info_i__max_slave__  = 0.025000000;
slave_timing[3][32+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][32+17].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+17].t_rxd1[0][1] = 2622ns;
slave_timing[3][32+17].t_rxd1[1][0] = 2774ns;
slave_timing[3][32+17].t_rxd1[0][2] = 1971ns;
slave_timing[3][32+17].t_rxd1[2][0] = 3332ns;
slave_timing[3][32+17].t_rxd2[0][2] = 3117ns;
slave_timing[3][32+17].t_rxd2[2][0] = 2175ns;
slave_timing[3][32+17].t_rxd2[1][2] = 2469ns;
slave_timing[3][32+17].t_rxd2[2][1] = 2966ns;

slave_timing[3][32+18].info_corner          = 2;
slave_timing[3][32+18].info_temp__j__       = 125;
slave_timing[3][32+18].info_i__quite_rec__  = 0.000000000;
slave_timing[3][32+18].info_dtr__ib__       = 1;
slave_timing[3][32+18].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+18].info_i__max_slave__  = 0.023000000;
slave_timing[3][32+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][32+18].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+18].t_rxd1[0][1] = 2792ns;
slave_timing[3][32+18].t_rxd1[1][0] = 2620ns;
slave_timing[3][32+18].t_rxd1[0][2] = 2061ns;
slave_timing[3][32+18].t_rxd1[2][0] = 3221ns;
slave_timing[3][32+18].t_rxd2[0][2] = 3473ns;
slave_timing[3][32+18].t_rxd2[2][0] = 1874ns;
slave_timing[3][32+18].t_rxd2[1][2] = 3053ns;
slave_timing[3][32+18].t_rxd2[2][1] = 2415ns;

slave_timing[3][32+19].info_corner          = 2;
slave_timing[3][32+19].info_temp__j__       = 125;
slave_timing[3][32+19].info_i__quite_rec__  = 0.000000000;
slave_timing[3][32+19].info_dtr__ib__       = 1;
slave_timing[3][32+19].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+19].info_i__max_slave__  = 0.025000000;
slave_timing[3][32+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][32+19].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+19].t_rxd1[0][1] = 2675ns;
slave_timing[3][32+19].t_rxd1[1][0] = 2703ns;
slave_timing[3][32+19].t_rxd1[0][2] = 1998ns;
slave_timing[3][32+19].t_rxd1[2][0] = 3276ns;
slave_timing[3][32+19].t_rxd2[0][2] = 3239ns;
slave_timing[3][32+19].t_rxd2[2][0] = 2046ns;
slave_timing[3][32+19].t_rxd2[1][2] = 2666ns;
slave_timing[3][32+19].t_rxd2[2][1] = 2694ns;

slave_timing[3][32+20].info_corner          = 2;
slave_timing[3][32+20].info_temp__j__       = 125;
slave_timing[3][32+20].info_i__quite_rec__  = 0.000000000;
slave_timing[3][32+20].info_dtr__ib__       = -1;
slave_timing[3][32+20].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+20].info_i__max_slave__  = 0.023000000;
slave_timing[3][32+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][32+20].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+20].t_rxd1[0][1] = 2912ns;
slave_timing[3][32+20].t_rxd1[1][0] = 2832ns;
slave_timing[3][32+20].t_rxd1[0][2] = 2202ns;
slave_timing[3][32+20].t_rxd1[2][0] = 3408ns;
slave_timing[3][32+20].t_rxd2[0][2] = 3328ns;
slave_timing[3][32+20].t_rxd2[2][0] = 2050ns;
slave_timing[3][32+20].t_rxd2[1][2] = 2775ns;
slave_timing[3][32+20].t_rxd2[2][1] = 2667ns;

slave_timing[3][32+21].info_corner          = 2;
slave_timing[3][32+21].info_temp__j__       = 125;
slave_timing[3][32+21].info_i__quite_rec__  = 0.000000000;
slave_timing[3][32+21].info_dtr__ib__       = -1;
slave_timing[3][32+21].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+21].info_i__max_slave__  = 0.025000000;
slave_timing[3][32+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][32+21].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+21].t_rxd1[0][1] = 2800ns;
slave_timing[3][32+21].t_rxd1[1][0] = 2905ns;
slave_timing[3][32+21].t_rxd1[0][2] = 2135ns;
slave_timing[3][32+21].t_rxd1[2][0] = 3459ns;
slave_timing[3][32+21].t_rxd2[0][2] = 3133ns;
slave_timing[3][32+21].t_rxd2[2][0] = 2196ns;
slave_timing[3][32+21].t_rxd2[1][2] = 2492ns;
slave_timing[3][32+21].t_rxd2[2][1] = 2944ns;

slave_timing[3][32+22].info_corner          = 2;
slave_timing[3][32+22].info_temp__j__       = 125;
slave_timing[3][32+22].info_i__quite_rec__  = 0.000000000;
slave_timing[3][32+22].info_dtr__ib__       = 1;
slave_timing[3][32+22].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+22].info_i__max_slave__  = 0.023000000;
slave_timing[3][32+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][32+22].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+22].t_rxd1[0][1] = 3021ns;
slave_timing[3][32+22].t_rxd1[1][0] = 2709ns;
slave_timing[3][32+22].t_rxd1[0][2] = 2224ns;
slave_timing[3][32+22].t_rxd1[2][0] = 3354ns;
slave_timing[3][32+22].t_rxd2[0][2] = 3488ns;
slave_timing[3][32+22].t_rxd2[2][0] = 1898ns;
slave_timing[3][32+22].t_rxd2[1][2] = 3066ns;
slave_timing[3][32+22].t_rxd2[2][1] = 2432ns;

slave_timing[3][32+23].info_corner          = 2;
slave_timing[3][32+23].info_temp__j__       = 125;
slave_timing[3][32+23].info_i__quite_rec__  = 0.000000000;
slave_timing[3][32+23].info_dtr__ib__       = 1;
slave_timing[3][32+23].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+23].info_i__max_slave__  = 0.025000000;
slave_timing[3][32+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][32+23].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+23].t_rxd1[0][1] = 2902ns;
slave_timing[3][32+23].t_rxd1[1][0] = 2841ns;
slave_timing[3][32+23].t_rxd1[0][2] = 2161ns;
slave_timing[3][32+23].t_rxd1[2][0] = 3409ns;
slave_timing[3][32+23].t_rxd2[0][2] = 3252ns;
slave_timing[3][32+23].t_rxd2[2][0] = 2070ns;
slave_timing[3][32+23].t_rxd2[1][2] = 2729ns;
slave_timing[3][32+23].t_rxd2[2][1] = 2714ns;

slave_timing[3][32+24].info_corner          = 2;
slave_timing[3][32+24].info_temp__j__       = 125;
slave_timing[3][32+24].info_i__quite_rec__  = 0.040000000;
slave_timing[3][32+24].info_dtr__ib__       = -1;
slave_timing[3][32+24].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+24].info_i__max_slave__  = 0.023000000;
slave_timing[3][32+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][32+24].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+24].t_rxd1[0][1] = 2746ns;
slave_timing[3][32+24].t_rxd1[1][0] = 2783ns;
slave_timing[3][32+24].t_rxd1[0][2] = 2058ns;
slave_timing[3][32+24].t_rxd1[2][0] = 3362ns;
slave_timing[3][32+24].t_rxd2[0][2] = 3510ns;
slave_timing[3][32+24].t_rxd2[2][0] = 2239ns;
slave_timing[3][32+24].t_rxd2[1][2] = 2938ns;
slave_timing[3][32+24].t_rxd2[2][1] = 2944ns;

slave_timing[3][32+25].info_corner          = 2;
slave_timing[3][32+25].info_temp__j__       = 125;
slave_timing[3][32+25].info_i__quite_rec__  = 0.040000000;
slave_timing[3][32+25].info_dtr__ib__       = -1;
slave_timing[3][32+25].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+25].info_i__max_slave__  = 0.025000000;
slave_timing[3][32+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][32+25].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+25].t_rxd1[0][1] = 2678ns;
slave_timing[3][32+25].t_rxd1[1][0] = 2828ns;
slave_timing[3][32+25].t_rxd1[0][2] = 1997ns;
slave_timing[3][32+25].t_rxd1[2][0] = 3408ns;
slave_timing[3][32+25].t_rxd2[0][2] = 3316ns;
slave_timing[3][32+25].t_rxd2[2][0] = 2384ns;
slave_timing[3][32+25].t_rxd2[1][2] = 2682ns;
slave_timing[3][32+25].t_rxd2[2][1] = 3200ns;

slave_timing[3][32+26].info_corner          = 2;
slave_timing[3][32+26].info_temp__j__       = 125;
slave_timing[3][32+26].info_i__quite_rec__  = 0.040000000;
slave_timing[3][32+26].info_dtr__ib__       = 1;
slave_timing[3][32+26].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+26].info_i__max_slave__  = 0.023000000;
slave_timing[3][32+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][32+26].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+26].t_rxd1[0][1] = 2853ns;
slave_timing[3][32+26].t_rxd1[1][0] = 2687ns;
slave_timing[3][32+26].t_rxd1[0][2] = 2122ns;
slave_timing[3][32+26].t_rxd1[2][0] = 3292ns;
slave_timing[3][32+26].t_rxd2[0][2] = 3714ns;
slave_timing[3][32+26].t_rxd2[2][0] = 2087ns;
slave_timing[3][32+26].t_rxd2[1][2] = 3226ns;
slave_timing[3][32+26].t_rxd2[2][1] = 2698ns;

slave_timing[3][32+27].info_corner          = 2;
slave_timing[3][32+27].info_temp__j__       = 125;
slave_timing[3][32+27].info_i__quite_rec__  = 0.040000000;
slave_timing[3][32+27].info_dtr__ib__       = 1;
slave_timing[3][32+27].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+27].info_i__max_slave__  = 0.025000000;
slave_timing[3][32+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][32+27].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+27].t_rxd1[0][1] = 2741ns;
slave_timing[3][32+27].t_rxd1[1][0] = 2772ns;
slave_timing[3][32+27].t_rxd1[0][2] = 2051ns;
slave_timing[3][32+27].t_rxd1[2][0] = 3350ns;
slave_timing[3][32+27].t_rxd2[0][2] = 3472ns;
slave_timing[3][32+27].t_rxd2[2][0] = 2259ns;
slave_timing[3][32+27].t_rxd2[1][2] = 2886ns;
slave_timing[3][32+27].t_rxd2[2][1] = 2989ns;

slave_timing[3][32+28].info_corner          = 2;
slave_timing[3][32+28].info_temp__j__       = 125;
slave_timing[3][32+28].info_i__quite_rec__  = 0.040000000;
slave_timing[3][32+28].info_dtr__ib__       = -1;
slave_timing[3][32+28].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+28].info_i__max_slave__  = 0.023000000;
slave_timing[3][32+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][32+28].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+28].t_rxd1[0][1] = 2798ns;
slave_timing[3][32+28].t_rxd1[1][0] = 2829ns;
slave_timing[3][32+28].t_rxd1[0][2] = 2133ns;
slave_timing[3][32+28].t_rxd1[2][0] = 3510ns;
slave_timing[3][32+28].t_rxd2[0][2] = 4066ns;
slave_timing[3][32+28].t_rxd2[2][0] = 2809ns;
slave_timing[3][32+28].t_rxd2[1][2] = 3555ns;
slave_timing[3][32+28].t_rxd2[2][1] = 3726ns;

slave_timing[3][32+29].info_corner          = 2;
slave_timing[3][32+29].info_temp__j__       = 125;
slave_timing[3][32+29].info_i__quite_rec__  = 0.040000000;
slave_timing[3][32+29].info_dtr__ib__       = -1;
slave_timing[3][32+29].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+29].info_i__max_slave__  = 0.025000000;
slave_timing[3][32+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][32+29].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+29].t_rxd1[0][1] = 2704ns;
slave_timing[3][32+29].t_rxd1[1][0] = 2907ns;
slave_timing[3][32+29].t_rxd1[0][2] = 2063ns;
slave_timing[3][32+29].t_rxd1[2][0] = 3636ns;
slave_timing[3][32+29].t_rxd2[0][2] = 3819ns;
slave_timing[3][32+29].t_rxd2[2][0] = 3004ns;
slave_timing[3][32+29].t_rxd2[1][2] = 3208ns;
slave_timing[3][32+29].t_rxd2[2][1] = 4085ns;

slave_timing[3][32+30].info_corner          = 2;
slave_timing[3][32+30].info_temp__j__       = 125;
slave_timing[3][32+30].info_i__quite_rec__  = 0.040000000;
slave_timing[3][32+30].info_dtr__ib__       = 1;
slave_timing[3][32+30].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+30].info_i__max_slave__  = 0.023000000;
slave_timing[3][32+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][32+30].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+30].t_rxd1[0][1] = 2911ns;
slave_timing[3][32+30].t_rxd1[1][0] = 2733ns;
slave_timing[3][32+30].t_rxd1[0][2] = 2185ns;
slave_timing[3][32+30].t_rxd1[2][0] = 3385ns;
slave_timing[3][32+30].t_rxd2[0][2] = 4333ns;
slave_timing[3][32+30].t_rxd2[2][0] = 2618ns;
slave_timing[3][32+30].t_rxd2[1][2] = 3894ns;
slave_timing[3][32+30].t_rxd2[2][1] = 3376ns;

slave_timing[3][32+31].info_corner          = 2;
slave_timing[3][32+31].info_temp__j__       = 125;
slave_timing[3][32+31].info_i__quite_rec__  = 0.040000000;
slave_timing[3][32+31].info_dtr__ib__       = 1;
slave_timing[3][32+31].info_i__offset_rec__ = 0.000000000;
slave_timing[3][32+31].info_i__max_slave__  = 0.025000000;
slave_timing[3][32+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][32+31].info_r__dsi_bus__    = 5.000;

slave_timing[3][32+31].t_rxd1[0][1] = 2796ns;
slave_timing[3][32+31].t_rxd1[1][0] = 2814ns;
slave_timing[3][32+31].t_rxd1[0][2] = 2121ns;
slave_timing[3][32+31].t_rxd1[2][0] = 3515ns;
slave_timing[3][32+31].t_rxd2[0][2] = 4011ns;
slave_timing[3][32+31].t_rxd2[2][0] = 2833ns;
slave_timing[3][32+31].t_rxd2[1][2] = 3485ns;
slave_timing[3][32+31].t_rxd2[2][1] = 3731ns;

//-----------------------------------------------------------------------------
// Copyright (c) 2023 Elmos SE
// Author     : Eugene - Easy UVM Generator
//
// Description: This file has been generated automatically by Eugene
//				This file should not be modified manually. 
//-----------------------------------------------------------------------------
`ifndef OSC_SEQUENCER_SV
`define OSC_SEQUENCER_SV

// You can insert code here by setting sequencer_inc_before_class in file osc.tpl

class osc_sequencer extends uvm_sequencer #(osc_tr);

	`uvm_component_utils(osc_sequencer)
	
	osc_config  m_config;

	function new(string name, uvm_component parent);
		super.new(name, parent);
	endfunction : new

	// You can insert code here by setting sequencer_inc_inside_class in file osc.tpl

endclass

typedef osc_sequencer osc_sequencer_t;

// You can insert code here by setting sequencer_inc_after_class in file osc.tpl

`endif



slave_timing[3][64+0].info_corner          = 3;
slave_timing[3][64+0].info_temp__j__       = 125;
slave_timing[3][64+0].info_i__quite_rec__  = 0.006000000;
slave_timing[3][64+0].info_dtr__ib__       = -1;
slave_timing[3][64+0].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+0].info_i__max_slave__  = 0.023000000;
slave_timing[3][64+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][64+0].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+0].t_rxd1[0][1] = 2748ns;
slave_timing[3][64+0].t_rxd1[1][0] = 2703ns;
slave_timing[3][64+0].t_rxd1[0][2] = 2031ns;
slave_timing[3][64+0].t_rxd1[2][0] = 3299ns;
slave_timing[3][64+0].t_rxd2[0][2] = 3287ns;
slave_timing[3][64+0].t_rxd2[2][0] = 2041ns;
slave_timing[3][64+0].t_rxd2[1][2] = 2748ns;
slave_timing[3][64+0].t_rxd2[2][1] = 2706ns;

slave_timing[3][64+1].info_corner          = 3;
slave_timing[3][64+1].info_temp__j__       = 125;
slave_timing[3][64+1].info_i__quite_rec__  = 0.006000000;
slave_timing[3][64+1].info_dtr__ib__       = -1;
slave_timing[3][64+1].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+1].info_i__max_slave__  = 0.025000000;
slave_timing[3][64+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][64+1].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+1].t_rxd1[0][1] = 2640ns;
slave_timing[3][64+1].t_rxd1[1][0] = 2784ns;
slave_timing[3][64+1].t_rxd1[0][2] = 1989ns;
slave_timing[3][64+1].t_rxd1[2][0] = 3350ns;
slave_timing[3][64+1].t_rxd2[0][2] = 3129ns;
slave_timing[3][64+1].t_rxd2[2][0] = 2190ns;
slave_timing[3][64+1].t_rxd2[1][2] = 2461ns;
slave_timing[3][64+1].t_rxd2[2][1] = 2989ns;

slave_timing[3][64+2].info_corner          = 3;
slave_timing[3][64+2].info_temp__j__       = 125;
slave_timing[3][64+2].info_i__quite_rec__  = 0.006000000;
slave_timing[3][64+2].info_dtr__ib__       = 1;
slave_timing[3][64+2].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+2].info_i__max_slave__  = 0.023000000;
slave_timing[3][64+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][64+2].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+2].t_rxd1[0][1] = 2809ns;
slave_timing[3][64+2].t_rxd1[1][0] = 2625ns;
slave_timing[3][64+2].t_rxd1[0][2] = 2072ns;
slave_timing[3][64+2].t_rxd1[2][0] = 3231ns;
slave_timing[3][64+2].t_rxd2[0][2] = 3480ns;
slave_timing[3][64+2].t_rxd2[2][0] = 1890ns;
slave_timing[3][64+2].t_rxd2[1][2] = 2983ns;
slave_timing[3][64+2].t_rxd2[2][1] = 2478ns;

slave_timing[3][64+3].info_corner          = 3;
slave_timing[3][64+3].info_temp__j__       = 125;
slave_timing[3][64+3].info_i__quite_rec__  = 0.006000000;
slave_timing[3][64+3].info_dtr__ib__       = 1;
slave_timing[3][64+3].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+3].info_i__max_slave__  = 0.025000000;
slave_timing[3][64+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][64+3].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+3].t_rxd1[0][1] = 2690ns;
slave_timing[3][64+3].t_rxd1[1][0] = 2703ns;
slave_timing[3][64+3].t_rxd1[0][2] = 2012ns;
slave_timing[3][64+3].t_rxd1[2][0] = 3288ns;
slave_timing[3][64+3].t_rxd2[0][2] = 3246ns;
slave_timing[3][64+3].t_rxd2[2][0] = 2066ns;
slave_timing[3][64+3].t_rxd2[1][2] = 2698ns;
slave_timing[3][64+3].t_rxd2[2][1] = 2723ns;

slave_timing[3][64+4].info_corner          = 3;
slave_timing[3][64+4].info_temp__j__       = 125;
slave_timing[3][64+4].info_i__quite_rec__  = 0.006000000;
slave_timing[3][64+4].info_dtr__ib__       = -1;
slave_timing[3][64+4].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+4].info_i__max_slave__  = 0.023000000;
slave_timing[3][64+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][64+4].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+4].t_rxd1[0][1] = 2944ns;
slave_timing[3][64+4].t_rxd1[1][0] = 2861ns;
slave_timing[3][64+4].t_rxd1[0][2] = 2225ns;
slave_timing[3][64+4].t_rxd1[2][0] = 3444ns;
slave_timing[3][64+4].t_rxd2[0][2] = 3344ns;
slave_timing[3][64+4].t_rxd2[2][0] = 2072ns;
slave_timing[3][64+4].t_rxd2[1][2] = 2778ns;
slave_timing[3][64+4].t_rxd2[2][1] = 2737ns;

slave_timing[3][64+5].info_corner          = 3;
slave_timing[3][64+5].info_temp__j__       = 125;
slave_timing[3][64+5].info_i__quite_rec__  = 0.006000000;
slave_timing[3][64+5].info_dtr__ib__       = -1;
slave_timing[3][64+5].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+5].info_i__max_slave__  = 0.025000000;
slave_timing[3][64+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][64+5].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+5].t_rxd1[0][1] = 2832ns;
slave_timing[3][64+5].t_rxd1[1][0] = 2940ns;
slave_timing[3][64+5].t_rxd1[0][2] = 2161ns;
slave_timing[3][64+5].t_rxd1[2][0] = 3497ns;
slave_timing[3][64+5].t_rxd2[0][2] = 3155ns;
slave_timing[3][64+5].t_rxd2[2][0] = 2217ns;
slave_timing[3][64+5].t_rxd2[1][2] = 2493ns;
slave_timing[3][64+5].t_rxd2[2][1] = 3016ns;

slave_timing[3][64+6].info_corner          = 3;
slave_timing[3][64+6].info_temp__j__       = 125;
slave_timing[3][64+6].info_i__quite_rec__  = 0.006000000;
slave_timing[3][64+6].info_dtr__ib__       = 1;
slave_timing[3][64+6].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+6].info_i__max_slave__  = 0.023000000;
slave_timing[3][64+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][64+6].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+6].t_rxd1[0][1] = 2991ns;
slave_timing[3][64+6].t_rxd1[1][0] = 2770ns;
slave_timing[3][64+6].t_rxd1[0][2] = 2237ns;
slave_timing[3][64+6].t_rxd1[2][0] = 3371ns;
slave_timing[3][64+6].t_rxd2[0][2] = 3499ns;
slave_timing[3][64+6].t_rxd2[2][0] = 1920ns;
slave_timing[3][64+6].t_rxd2[1][2] = 3058ns;
slave_timing[3][64+6].t_rxd2[2][1] = 2469ns;

slave_timing[3][64+7].info_corner          = 3;
slave_timing[3][64+7].info_temp__j__       = 125;
slave_timing[3][64+7].info_i__quite_rec__  = 0.006000000;
slave_timing[3][64+7].info_dtr__ib__       = 1;
slave_timing[3][64+7].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+7].info_i__max_slave__  = 0.025000000;
slave_timing[3][64+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][64+7].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+7].t_rxd1[0][1] = 2874ns;
slave_timing[3][64+7].t_rxd1[1][0] = 2852ns;
slave_timing[3][64+7].t_rxd1[0][2] = 2175ns;
slave_timing[3][64+7].t_rxd1[2][0] = 3426ns;
slave_timing[3][64+7].t_rxd2[0][2] = 3275ns;
slave_timing[3][64+7].t_rxd2[2][0] = 2095ns;
slave_timing[3][64+7].t_rxd2[1][2] = 2721ns;
slave_timing[3][64+7].t_rxd2[2][1] = 2750ns;

slave_timing[3][64+8].info_corner          = 3;
slave_timing[3][64+8].info_temp__j__       = 125;
slave_timing[3][64+8].info_i__quite_rec__  = 0.003000000;
slave_timing[3][64+8].info_dtr__ib__       = -1;
slave_timing[3][64+8].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+8].info_i__max_slave__  = 0.023000000;
slave_timing[3][64+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][64+8].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+8].t_rxd1[0][1] = 2680ns;
slave_timing[3][64+8].t_rxd1[1][0] = 2700ns;
slave_timing[3][64+8].t_rxd1[0][2] = 2007ns;
slave_timing[3][64+8].t_rxd1[2][0] = 3277ns;
slave_timing[3][64+8].t_rxd2[0][2] = 3271ns;
slave_timing[3][64+8].t_rxd2[2][0] = 2024ns;
slave_timing[3][64+8].t_rxd2[1][2] = 2710ns;
slave_timing[3][64+8].t_rxd2[2][1] = 2691ns;

slave_timing[3][64+9].info_corner          = 3;
slave_timing[3][64+9].info_temp__j__       = 125;
slave_timing[3][64+9].info_i__quite_rec__  = 0.003000000;
slave_timing[3][64+9].info_dtr__ib__       = -1;
slave_timing[3][64+9].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+9].info_i__max_slave__  = 0.025000000;
slave_timing[3][64+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][64+9].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+9].t_rxd1[0][1] = 2583ns;
slave_timing[3][64+9].t_rxd1[1][0] = 2780ns;
slave_timing[3][64+9].t_rxd1[0][2] = 1920ns;
slave_timing[3][64+9].t_rxd1[2][0] = 3331ns;
slave_timing[3][64+9].t_rxd2[0][2] = 3058ns;
slave_timing[3][64+9].t_rxd2[2][0] = 2170ns;
slave_timing[3][64+9].t_rxd2[1][2] = 2427ns;
slave_timing[3][64+9].t_rxd2[2][1] = 2970ns;

slave_timing[3][64+10].info_corner          = 3;
slave_timing[3][64+10].info_temp__j__       = 125;
slave_timing[3][64+10].info_i__quite_rec__  = 0.003000000;
slave_timing[3][64+10].info_dtr__ib__       = 1;
slave_timing[3][64+10].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+10].info_i__max_slave__  = 0.023000000;
slave_timing[3][64+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][64+10].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+10].t_rxd1[0][1] = 2779ns;
slave_timing[3][64+10].t_rxd1[1][0] = 2575ns;
slave_timing[3][64+10].t_rxd1[0][2] = 2053ns;
slave_timing[3][64+10].t_rxd1[2][0] = 3185ns;
slave_timing[3][64+10].t_rxd2[0][2] = 3462ns;
slave_timing[3][64+10].t_rxd2[2][0] = 1855ns;
slave_timing[3][64+10].t_rxd2[1][2] = 2984ns;
slave_timing[3][64+10].t_rxd2[2][1] = 2426ns;

slave_timing[3][64+11].info_corner          = 3;
slave_timing[3][64+11].info_temp__j__       = 125;
slave_timing[3][64+11].info_i__quite_rec__  = 0.003000000;
slave_timing[3][64+11].info_dtr__ib__       = 1;
slave_timing[3][64+11].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+11].info_i__max_slave__  = 0.025000000;
slave_timing[3][64+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][64+11].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+11].t_rxd1[0][1] = 2664ns;
slave_timing[3][64+11].t_rxd1[1][0] = 2657ns;
slave_timing[3][64+11].t_rxd1[0][2] = 1984ns;
slave_timing[3][64+11].t_rxd1[2][0] = 3240ns;
slave_timing[3][64+11].t_rxd2[0][2] = 3228ns;
slave_timing[3][64+11].t_rxd2[2][0] = 2030ns;
slave_timing[3][64+11].t_rxd2[1][2] = 2653ns;
slave_timing[3][64+11].t_rxd2[2][1] = 2707ns;

slave_timing[3][64+12].info_corner          = 3;
slave_timing[3][64+12].info_temp__j__       = 125;
slave_timing[3][64+12].info_i__quite_rec__  = 0.003000000;
slave_timing[3][64+12].info_dtr__ib__       = -1;
slave_timing[3][64+12].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+12].info_i__max_slave__  = 0.023000000;
slave_timing[3][64+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][64+12].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+12].t_rxd1[0][1] = 2933ns;
slave_timing[3][64+12].t_rxd1[1][0] = 2825ns;
slave_timing[3][64+12].t_rxd1[0][2] = 2194ns;
slave_timing[3][64+12].t_rxd1[2][0] = 3437ns;
slave_timing[3][64+12].t_rxd2[0][2] = 3301ns;
slave_timing[3][64+12].t_rxd2[2][0] = 2055ns;
slave_timing[3][64+12].t_rxd2[1][2] = 2775ns;
slave_timing[3][64+12].t_rxd2[2][1] = 2681ns;

slave_timing[3][64+13].info_corner          = 3;
slave_timing[3][64+13].info_temp__j__       = 125;
slave_timing[3][64+13].info_i__quite_rec__  = 0.003000000;
slave_timing[3][64+13].info_dtr__ib__       = -1;
slave_timing[3][64+13].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+13].info_i__max_slave__  = 0.025000000;
slave_timing[3][64+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][64+13].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+13].t_rxd1[0][1] = 2824ns;
slave_timing[3][64+13].t_rxd1[1][0] = 2903ns;
slave_timing[3][64+13].t_rxd1[0][2] = 2129ns;
slave_timing[3][64+13].t_rxd1[2][0] = 3488ns;
slave_timing[3][64+13].t_rxd2[0][2] = 3111ns;
slave_timing[3][64+13].t_rxd2[2][0] = 2201ns;
slave_timing[3][64+13].t_rxd2[1][2] = 2487ns;
slave_timing[3][64+13].t_rxd2[2][1] = 2959ns;

slave_timing[3][64+14].info_corner          = 3;
slave_timing[3][64+14].info_temp__j__       = 125;
slave_timing[3][64+14].info_i__quite_rec__  = 0.003000000;
slave_timing[3][64+14].info_dtr__ib__       = 1;
slave_timing[3][64+14].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+14].info_i__max_slave__  = 0.023000000;
slave_timing[3][64+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][64+14].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+14].t_rxd1[0][1] = 2976ns;
slave_timing[3][64+14].t_rxd1[1][0] = 2727ns;
slave_timing[3][64+14].t_rxd1[0][2] = 2229ns;
slave_timing[3][64+14].t_rxd1[2][0] = 3326ns;
slave_timing[3][64+14].t_rxd2[0][2] = 3485ns;
slave_timing[3][64+14].t_rxd2[2][0] = 1881ns;
slave_timing[3][64+14].t_rxd2[1][2] = 3008ns;
slave_timing[3][64+14].t_rxd2[2][1] = 2455ns;

slave_timing[3][64+15].info_corner          = 3;
slave_timing[3][64+15].info_temp__j__       = 125;
slave_timing[3][64+15].info_i__quite_rec__  = 0.003000000;
slave_timing[3][64+15].info_dtr__ib__       = 1;
slave_timing[3][64+15].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+15].info_i__max_slave__  = 0.025000000;
slave_timing[3][64+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][64+15].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+15].t_rxd1[0][1] = 2859ns;
slave_timing[3][64+15].t_rxd1[1][0] = 2808ns;
slave_timing[3][64+15].t_rxd1[0][2] = 2163ns;
slave_timing[3][64+15].t_rxd1[2][0] = 3381ns;
slave_timing[3][64+15].t_rxd2[0][2] = 3253ns;
slave_timing[3][64+15].t_rxd2[2][0] = 2050ns;
slave_timing[3][64+15].t_rxd2[1][2] = 2683ns;
slave_timing[3][64+15].t_rxd2[2][1] = 2733ns;

slave_timing[3][64+16].info_corner          = 3;
slave_timing[3][64+16].info_temp__j__       = 125;
slave_timing[3][64+16].info_i__quite_rec__  = 0.000000000;
slave_timing[3][64+16].info_dtr__ib__       = -1;
slave_timing[3][64+16].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+16].info_i__max_slave__  = 0.023000000;
slave_timing[3][64+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][64+16].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+16].t_rxd1[0][1] = 2674ns;
slave_timing[3][64+16].t_rxd1[1][0] = 2657ns;
slave_timing[3][64+16].t_rxd1[0][2] = 1991ns;
slave_timing[3][64+16].t_rxd1[2][0] = 3232ns;
slave_timing[3][64+16].t_rxd2[0][2] = 3248ns;
slave_timing[3][64+16].t_rxd2[2][0] = 1988ns;
slave_timing[3][64+16].t_rxd2[1][2] = 2696ns;
slave_timing[3][64+16].t_rxd2[2][1] = 2649ns;

slave_timing[3][64+17].info_corner          = 3;
slave_timing[3][64+17].info_temp__j__       = 125;
slave_timing[3][64+17].info_i__quite_rec__  = 0.000000000;
slave_timing[3][64+17].info_dtr__ib__       = -1;
slave_timing[3][64+17].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+17].info_i__max_slave__  = 0.025000000;
slave_timing[3][64+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][64+17].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+17].t_rxd1[0][1] = 2572ns;
slave_timing[3][64+17].t_rxd1[1][0] = 2733ns;
slave_timing[3][64+17].t_rxd1[0][2] = 1926ns;
slave_timing[3][64+17].t_rxd1[2][0] = 3280ns;
slave_timing[3][64+17].t_rxd2[0][2] = 3050ns;
slave_timing[3][64+17].t_rxd2[2][0] = 2138ns;
slave_timing[3][64+17].t_rxd2[1][2] = 2411ns;
slave_timing[3][64+17].t_rxd2[2][1] = 2921ns;

slave_timing[3][64+18].info_corner          = 3;
slave_timing[3][64+18].info_temp__j__       = 125;
slave_timing[3][64+18].info_i__quite_rec__  = 0.000000000;
slave_timing[3][64+18].info_dtr__ib__       = 1;
slave_timing[3][64+18].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+18].info_i__max_slave__  = 0.023000000;
slave_timing[3][64+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][64+18].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+18].t_rxd1[0][1] = 2770ns;
slave_timing[3][64+18].t_rxd1[1][0] = 2539ns;
slave_timing[3][64+18].t_rxd1[0][2] = 2042ns;
slave_timing[3][64+18].t_rxd1[2][0] = 3146ns;
slave_timing[3][64+18].t_rxd2[0][2] = 3433ns;
slave_timing[3][64+18].t_rxd2[2][0] = 1817ns;
slave_timing[3][64+18].t_rxd2[1][2] = 3012ns;
slave_timing[3][64+18].t_rxd2[2][1] = 2345ns;

slave_timing[3][64+19].info_corner          = 3;
slave_timing[3][64+19].info_temp__j__       = 125;
slave_timing[3][64+19].info_i__quite_rec__  = 0.000000000;
slave_timing[3][64+19].info_dtr__ib__       = 1;
slave_timing[3][64+19].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+19].info_i__max_slave__  = 0.025000000;
slave_timing[3][64+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][64+19].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+19].t_rxd1[0][1] = 2651ns;
slave_timing[3][64+19].t_rxd1[1][0] = 2624ns;
slave_timing[3][64+19].t_rxd1[0][2] = 1977ns;
slave_timing[3][64+19].t_rxd1[2][0] = 3199ns;
slave_timing[3][64+19].t_rxd2[0][2] = 3199ns;
slave_timing[3][64+19].t_rxd2[2][0] = 1993ns;
slave_timing[3][64+19].t_rxd2[1][2] = 2636ns;
slave_timing[3][64+19].t_rxd2[2][1] = 2661ns;

slave_timing[3][64+20].info_corner          = 3;
slave_timing[3][64+20].info_temp__j__       = 125;
slave_timing[3][64+20].info_i__quite_rec__  = 0.000000000;
slave_timing[3][64+20].info_dtr__ib__       = -1;
slave_timing[3][64+20].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+20].info_i__max_slave__  = 0.023000000;
slave_timing[3][64+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][64+20].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+20].t_rxd1[0][1] = 2898ns;
slave_timing[3][64+20].t_rxd1[1][0] = 2813ns;
slave_timing[3][64+20].t_rxd1[0][2] = 2195ns;
slave_timing[3][64+20].t_rxd1[2][0] = 3376ns;
slave_timing[3][64+20].t_rxd2[0][2] = 3268ns;
slave_timing[3][64+20].t_rxd2[2][0] = 2018ns;
slave_timing[3][64+20].t_rxd2[1][2] = 2714ns;
slave_timing[3][64+20].t_rxd2[2][1] = 2667ns;

slave_timing[3][64+21].info_corner          = 3;
slave_timing[3][64+21].info_temp__j__       = 125;
slave_timing[3][64+21].info_i__quite_rec__  = 0.000000000;
slave_timing[3][64+21].info_dtr__ib__       = -1;
slave_timing[3][64+21].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+21].info_i__max_slave__  = 0.025000000;
slave_timing[3][64+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][64+21].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+21].t_rxd1[0][1] = 2793ns;
slave_timing[3][64+21].t_rxd1[1][0] = 2891ns;
slave_timing[3][64+21].t_rxd1[0][2] = 2133ns;
slave_timing[3][64+21].t_rxd1[2][0] = 3429ns;
slave_timing[3][64+21].t_rxd2[0][2] = 3077ns;
slave_timing[3][64+21].t_rxd2[2][0] = 2166ns;
slave_timing[3][64+21].t_rxd2[1][2] = 2434ns;
slave_timing[3][64+21].t_rxd2[2][1] = 2910ns;

slave_timing[3][64+22].info_corner          = 3;
slave_timing[3][64+22].info_temp__j__       = 125;
slave_timing[3][64+22].info_i__quite_rec__  = 0.000000000;
slave_timing[3][64+22].info_dtr__ib__       = 1;
slave_timing[3][64+22].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+22].info_i__max_slave__  = 0.023000000;
slave_timing[3][64+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][64+22].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+22].t_rxd1[0][1] = 2985ns;
slave_timing[3][64+22].t_rxd1[1][0] = 2691ns;
slave_timing[3][64+22].t_rxd1[0][2] = 2232ns;
slave_timing[3][64+22].t_rxd1[2][0] = 3284ns;
slave_timing[3][64+22].t_rxd2[0][2] = 3453ns;
slave_timing[3][64+22].t_rxd2[2][0] = 1842ns;
slave_timing[3][64+22].t_rxd2[1][2] = 3037ns;
slave_timing[3][64+22].t_rxd2[2][1] = 2370ns;

slave_timing[3][64+23].info_corner          = 3;
slave_timing[3][64+23].info_temp__j__       = 125;
slave_timing[3][64+23].info_i__quite_rec__  = 0.000000000;
slave_timing[3][64+23].info_dtr__ib__       = 1;
slave_timing[3][64+23].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+23].info_i__max_slave__  = 0.025000000;
slave_timing[3][64+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][64+23].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+23].t_rxd1[0][1] = 2868ns;
slave_timing[3][64+23].t_rxd1[1][0] = 2773ns;
slave_timing[3][64+23].t_rxd1[0][2] = 2167ns;
slave_timing[3][64+23].t_rxd1[2][0] = 3337ns;
slave_timing[3][64+23].t_rxd2[0][2] = 3220ns;
slave_timing[3][64+23].t_rxd2[2][0] = 2014ns;
slave_timing[3][64+23].t_rxd2[1][2] = 2662ns;
slave_timing[3][64+23].t_rxd2[2][1] = 2683ns;

slave_timing[3][64+24].info_corner          = 3;
slave_timing[3][64+24].info_temp__j__       = 125;
slave_timing[3][64+24].info_i__quite_rec__  = 0.040000000;
slave_timing[3][64+24].info_dtr__ib__       = -1;
slave_timing[3][64+24].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+24].info_i__max_slave__  = 0.023000000;
slave_timing[3][64+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][64+24].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+24].t_rxd1[0][1] = 2759ns;
slave_timing[3][64+24].t_rxd1[1][0] = 2760ns;
slave_timing[3][64+24].t_rxd1[0][2] = 2067ns;
slave_timing[3][64+24].t_rxd1[2][0] = 3350ns;
slave_timing[3][64+24].t_rxd2[0][2] = 3332ns;
slave_timing[3][64+24].t_rxd2[2][0] = 2046ns;
slave_timing[3][64+24].t_rxd2[1][2] = 2741ns;
slave_timing[3][64+24].t_rxd2[2][1] = 2707ns;

slave_timing[3][64+25].info_corner          = 3;
slave_timing[3][64+25].info_temp__j__       = 125;
slave_timing[3][64+25].info_i__quite_rec__  = 0.040000000;
slave_timing[3][64+25].info_dtr__ib__       = -1;
slave_timing[3][64+25].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+25].info_i__max_slave__  = 0.025000000;
slave_timing[3][64+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][64+25].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+25].t_rxd1[0][1] = 2653ns;
slave_timing[3][64+25].t_rxd1[1][0] = 2842ns;
slave_timing[3][64+25].t_rxd1[0][2] = 2004ns;
slave_timing[3][64+25].t_rxd1[2][0] = 3401ns;
slave_timing[3][64+25].t_rxd2[0][2] = 3148ns;
slave_timing[3][64+25].t_rxd2[2][0] = 2200ns;
slave_timing[3][64+25].t_rxd2[1][2] = 2460ns;
slave_timing[3][64+25].t_rxd2[2][1] = 2989ns;

slave_timing[3][64+26].info_corner          = 3;
slave_timing[3][64+26].info_temp__j__       = 125;
slave_timing[3][64+26].info_i__quite_rec__  = 0.040000000;
slave_timing[3][64+26].info_dtr__ib__       = 1;
slave_timing[3][64+26].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+26].info_i__max_slave__  = 0.023000000;
slave_timing[3][64+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][64+26].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+26].t_rxd1[0][1] = 2835ns;
slave_timing[3][64+26].t_rxd1[1][0] = 2693ns;
slave_timing[3][64+26].t_rxd1[0][2] = 2110ns;
slave_timing[3][64+26].t_rxd1[2][0] = 3305ns;
slave_timing[3][64+26].t_rxd2[0][2] = 3501ns;
slave_timing[3][64+26].t_rxd2[2][0] = 1920ns;
slave_timing[3][64+26].t_rxd2[1][2] = 2983ns;
slave_timing[3][64+26].t_rxd2[2][1] = 2508ns;

slave_timing[3][64+27].info_corner          = 3;
slave_timing[3][64+27].info_temp__j__       = 125;
slave_timing[3][64+27].info_i__quite_rec__  = 0.040000000;
slave_timing[3][64+27].info_dtr__ib__       = 1;
slave_timing[3][64+27].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+27].info_i__max_slave__  = 0.025000000;
slave_timing[3][64+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][64+27].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+27].t_rxd1[0][1] = 2724ns;
slave_timing[3][64+27].t_rxd1[1][0] = 2777ns;
slave_timing[3][64+27].t_rxd1[0][2] = 2021ns;
slave_timing[3][64+27].t_rxd1[2][0] = 3358ns;
slave_timing[3][64+27].t_rxd2[0][2] = 3258ns;
slave_timing[3][64+27].t_rxd2[2][0] = 2105ns;
slave_timing[3][64+27].t_rxd2[1][2] = 2665ns;
slave_timing[3][64+27].t_rxd2[2][1] = 2795ns;

slave_timing[3][64+28].info_corner          = 3;
slave_timing[3][64+28].info_temp__j__       = 125;
slave_timing[3][64+28].info_i__quite_rec__  = 0.040000000;
slave_timing[3][64+28].info_dtr__ib__       = -1;
slave_timing[3][64+28].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+28].info_i__max_slave__  = 0.023000000;
slave_timing[3][64+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][64+28].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+28].t_rxd1[0][1] = 2849ns;
slave_timing[3][64+28].t_rxd1[1][0] = 2845ns;
slave_timing[3][64+28].t_rxd1[0][2] = 2158ns;
slave_timing[3][64+28].t_rxd1[2][0] = 3386ns;
slave_timing[3][64+28].t_rxd2[0][2] = 3391ns;
slave_timing[3][64+28].t_rxd2[2][0] = 2350ns;
slave_timing[3][64+28].t_rxd2[1][2] = 2809ns;
slave_timing[3][64+28].t_rxd2[2][1] = 2971ns;

slave_timing[3][64+29].info_corner          = 3;
slave_timing[3][64+29].info_temp__j__       = 125;
slave_timing[3][64+29].info_i__quite_rec__  = 0.040000000;
slave_timing[3][64+29].info_dtr__ib__       = -1;
slave_timing[3][64+29].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+29].info_i__max_slave__  = 0.025000000;
slave_timing[3][64+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][64+29].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+29].t_rxd1[0][1] = 2746ns;
slave_timing[3][64+29].t_rxd1[1][0] = 2922ns;
slave_timing[3][64+29].t_rxd1[0][2] = 2094ns;
slave_timing[3][64+29].t_rxd1[2][0] = 3390ns;
slave_timing[3][64+29].t_rxd2[0][2] = 3216ns;
slave_timing[3][64+29].t_rxd2[2][0] = 2568ns;
slave_timing[3][64+29].t_rxd2[1][2] = 2526ns;
slave_timing[3][64+29].t_rxd2[2][1] = 3334ns;

slave_timing[3][64+30].info_corner          = 3;
slave_timing[3][64+30].info_temp__j__       = 125;
slave_timing[3][64+30].info_i__quite_rec__  = 0.040000000;
slave_timing[3][64+30].info_dtr__ib__       = 1;
slave_timing[3][64+30].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+30].info_i__max_slave__  = 0.023000000;
slave_timing[3][64+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][64+30].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+30].t_rxd1[0][1] = 2923ns;
slave_timing[3][64+30].t_rxd1[1][0] = 2775ns;
slave_timing[3][64+30].t_rxd1[0][2] = 2194ns;
slave_timing[3][64+30].t_rxd1[2][0] = 3357ns;
slave_timing[3][64+30].t_rxd2[0][2] = 3565ns;
slave_timing[3][64+30].t_rxd2[2][0] = 2216ns;
slave_timing[3][64+30].t_rxd2[1][2] = 3046ns;
slave_timing[3][64+30].t_rxd2[2][1] = 2761ns;

slave_timing[3][64+31].info_corner          = 3;
slave_timing[3][64+31].info_temp__j__       = 125;
slave_timing[3][64+31].info_i__quite_rec__  = 0.040000000;
slave_timing[3][64+31].info_dtr__ib__       = 1;
slave_timing[3][64+31].info_i__offset_rec__ = 0.000000000;
slave_timing[3][64+31].info_i__max_slave__  = 0.025000000;
slave_timing[3][64+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][64+31].info_r__dsi_bus__    = 5.000;

slave_timing[3][64+31].t_rxd1[0][1] = 2808ns;
slave_timing[3][64+31].t_rxd1[1][0] = 2860ns;
slave_timing[3][64+31].t_rxd1[0][2] = 2131ns;
slave_timing[3][64+31].t_rxd1[2][0] = 3380ns;
slave_timing[3][64+31].t_rxd2[0][2] = 3358ns;
slave_timing[3][64+31].t_rxd2[2][0] = 2451ns;
slave_timing[3][64+31].t_rxd2[1][2] = 2736ns;
slave_timing[3][64+31].t_rxd2[2][1] = 3144ns;

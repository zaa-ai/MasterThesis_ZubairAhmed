
slave_timing[0][0].info_corner          = 1;
slave_timing[0][0].info_temp__j__       = 125;
slave_timing[0][0].info_i__quite_rec__  = 0.006000000;
slave_timing[0][0].info_dtr__ib__       = -1;
slave_timing[0][0].info_i__offset_rec__ = 0.000000000;
slave_timing[0][0].info_i__max_slave__  = 0.023000000;
slave_timing[0][0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][0].info_r__dsi_bus__    = 5.000;

slave_timing[0][0].t_rxd1[0][1] = 1098ns;
slave_timing[0][0].t_rxd1[1][0] = 1111ns;
slave_timing[0][0].t_rxd1[0][2] = 818ns;
slave_timing[0][0].t_rxd1[2][0] = 1364ns;
slave_timing[0][0].t_rxd2[0][2] = 1320ns;
slave_timing[0][0].t_rxd2[2][0] = 815ns;
slave_timing[0][0].t_rxd2[1][2] = 1067ns;
slave_timing[0][0].t_rxd2[2][1] = 1080ns;

slave_timing[0][1].info_corner          = 1;
slave_timing[0][1].info_temp__j__       = 125;
slave_timing[0][1].info_i__quite_rec__  = 0.006000000;
slave_timing[0][1].info_dtr__ib__       = -1;
slave_timing[0][1].info_i__offset_rec__ = 0.000000000;
slave_timing[0][1].info_i__max_slave__  = 0.025000000;
slave_timing[0][1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][1].info_r__dsi_bus__    = 5.000;

slave_timing[0][1].t_rxd1[0][1] = 1052ns;
slave_timing[0][1].t_rxd1[1][0] = 1143ns;
slave_timing[0][1].t_rxd1[0][2] = 795ns;
slave_timing[0][1].t_rxd1[2][0] = 1390ns;
slave_timing[0][1].t_rxd2[0][2] = 1228ns;
slave_timing[0][1].t_rxd2[2][0] = 864ns;
slave_timing[0][1].t_rxd2[1][2] = 949ns;
slave_timing[0][1].t_rxd2[2][1] = 1200ns;

slave_timing[0][2].info_corner          = 1;
slave_timing[0][2].info_temp__j__       = 125;
slave_timing[0][2].info_i__quite_rec__  = 0.006000000;
slave_timing[0][2].info_dtr__ib__       = 1;
slave_timing[0][2].info_i__offset_rec__ = 0.000000000;
slave_timing[0][2].info_i__max_slave__  = 0.023000000;
slave_timing[0][2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][2].info_r__dsi_bus__    = 5.000;

slave_timing[0][2].t_rxd1[0][1] = 1134ns;
slave_timing[0][2].t_rxd1[1][0] = 1064ns;
slave_timing[0][2].t_rxd1[0][2] = 833ns;
slave_timing[0][2].t_rxd1[2][0] = 1323ns;
slave_timing[0][2].t_rxd2[0][2] = 1422ns;
slave_timing[0][2].t_rxd2[2][0] = 761ns;
slave_timing[0][2].t_rxd2[1][2] = 1191ns;
slave_timing[0][2].t_rxd2[2][1] = 976ns;

slave_timing[0][3].info_corner          = 1;
slave_timing[0][3].info_temp__j__       = 125;
slave_timing[0][3].info_i__quite_rec__  = 0.006000000;
slave_timing[0][3].info_dtr__ib__       = 1;
slave_timing[0][3].info_i__offset_rec__ = 0.000000000;
slave_timing[0][3].info_i__max_slave__  = 0.025000000;
slave_timing[0][3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][3].info_r__dsi_bus__    = 5.000;

slave_timing[0][3].t_rxd1[0][1] = 1084ns;
slave_timing[0][3].t_rxd1[1][0] = 1101ns;
slave_timing[0][3].t_rxd1[0][2] = 807ns;
slave_timing[0][3].t_rxd1[2][0] = 1350ns;
slave_timing[0][3].t_rxd2[0][2] = 1298ns;
slave_timing[0][3].t_rxd2[2][0] = 816ns;
slave_timing[0][3].t_rxd2[1][2] = 1049ns;
slave_timing[0][3].t_rxd2[2][1] = 1092ns;

slave_timing[0][4].info_corner          = 1;
slave_timing[0][4].info_temp__j__       = 125;
slave_timing[0][4].info_i__quite_rec__  = 0.006000000;
slave_timing[0][4].info_dtr__ib__       = -1;
slave_timing[0][4].info_i__offset_rec__ = 0.000000000;
slave_timing[0][4].info_i__max_slave__  = 0.023000000;
slave_timing[0][4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][4].info_r__dsi_bus__    = 5.000;

slave_timing[0][4].t_rxd1[0][1] = 1293ns;
slave_timing[0][4].t_rxd1[1][0] = 1262ns;
slave_timing[0][4].t_rxd1[0][2] = 960ns;
slave_timing[0][4].t_rxd1[2][0] = 1504ns;
slave_timing[0][4].t_rxd2[0][2] = 1382ns;
slave_timing[0][4].t_rxd2[2][0] = 854ns;
slave_timing[0][4].t_rxd2[1][2] = 1095ns;
slave_timing[0][4].t_rxd2[2][1] = 1110ns;

slave_timing[0][5].info_corner          = 1;
slave_timing[0][5].info_temp__j__       = 125;
slave_timing[0][5].info_i__quite_rec__  = 0.006000000;
slave_timing[0][5].info_dtr__ib__       = -1;
slave_timing[0][5].info_i__offset_rec__ = 0.000000000;
slave_timing[0][5].info_i__max_slave__  = 0.025000000;
slave_timing[0][5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][5].info_r__dsi_bus__    = 5.000;

slave_timing[0][5].t_rxd1[0][1] = 1239ns;
slave_timing[0][5].t_rxd1[1][0] = 1294ns;
slave_timing[0][5].t_rxd1[0][2] = 933ns;
slave_timing[0][5].t_rxd1[2][0] = 1529ns;
slave_timing[0][5].t_rxd2[0][2] = 1290ns;
slave_timing[0][5].t_rxd2[2][0] = 905ns;
slave_timing[0][5].t_rxd2[1][2] = 982ns;
slave_timing[0][5].t_rxd2[2][1] = 1224ns;

slave_timing[0][6].info_corner          = 1;
slave_timing[0][6].info_temp__j__       = 125;
slave_timing[0][6].info_i__quite_rec__  = 0.006000000;
slave_timing[0][6].info_dtr__ib__       = 1;
slave_timing[0][6].info_i__offset_rec__ = 0.000000000;
slave_timing[0][6].info_i__max_slave__  = 0.023000000;
slave_timing[0][6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][6].info_r__dsi_bus__    = 5.000;

slave_timing[0][6].t_rxd1[0][1] = 1342ns;
slave_timing[0][6].t_rxd1[1][0] = 1211ns;
slave_timing[0][6].t_rxd1[0][2] = 977ns;
slave_timing[0][6].t_rxd1[2][0] = 1462ns;
slave_timing[0][6].t_rxd2[0][2] = 1483ns;
slave_timing[0][6].t_rxd2[2][0] = 798ns;
slave_timing[0][6].t_rxd2[1][2] = 1215ns;
slave_timing[0][6].t_rxd2[2][1] = 1010ns;

slave_timing[0][7].info_corner          = 1;
slave_timing[0][7].info_temp__j__       = 125;
slave_timing[0][7].info_i__quite_rec__  = 0.006000000;
slave_timing[0][7].info_dtr__ib__       = 1;
slave_timing[0][7].info_i__offset_rec__ = 0.000000000;
slave_timing[0][7].info_i__max_slave__  = 0.025000000;
slave_timing[0][7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][7].info_r__dsi_bus__    = 5.000;

slave_timing[0][7].t_rxd1[0][1] = 1278ns;
slave_timing[0][7].t_rxd1[1][0] = 1245ns;
slave_timing[0][7].t_rxd1[0][2] = 948ns;
slave_timing[0][7].t_rxd1[2][0] = 1489ns;
slave_timing[0][7].t_rxd2[0][2] = 1361ns;
slave_timing[0][7].t_rxd2[2][0] = 857ns;
slave_timing[0][7].t_rxd2[1][2] = 1076ns;
slave_timing[0][7].t_rxd2[2][1] = 1117ns;

slave_timing[0][8].info_corner          = 1;
slave_timing[0][8].info_temp__j__       = 125;
slave_timing[0][8].info_i__quite_rec__  = 0.003000000;
slave_timing[0][8].info_dtr__ib__       = -1;
slave_timing[0][8].info_i__offset_rec__ = 0.000000000;
slave_timing[0][8].info_i__max_slave__  = 0.023000000;
slave_timing[0][8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][8].info_r__dsi_bus__    = 5.000;

slave_timing[0][8].t_rxd1[0][1] = 1075ns;
slave_timing[0][8].t_rxd1[1][0] = 1104ns;
slave_timing[0][8].t_rxd1[0][2] = 805ns;
slave_timing[0][8].t_rxd1[2][0] = 1352ns;
slave_timing[0][8].t_rxd2[0][2] = 1301ns;
slave_timing[0][8].t_rxd2[2][0] = 816ns;
slave_timing[0][8].t_rxd2[1][2] = 1051ns;
slave_timing[0][8].t_rxd2[2][1] = 1086ns;

slave_timing[0][9].info_corner          = 1;
slave_timing[0][9].info_temp__j__       = 125;
slave_timing[0][9].info_i__quite_rec__  = 0.003000000;
slave_timing[0][9].info_dtr__ib__       = -1;
slave_timing[0][9].info_i__offset_rec__ = 0.000000000;
slave_timing[0][9].info_i__max_slave__  = 0.025000000;
slave_timing[0][9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][9].info_r__dsi_bus__    = 5.000;

slave_timing[0][9].t_rxd1[0][1] = 1029ns;
slave_timing[0][9].t_rxd1[1][0] = 1135ns;
slave_timing[0][9].t_rxd1[0][2] = 779ns;
slave_timing[0][9].t_rxd1[2][0] = 1376ns;
slave_timing[0][9].t_rxd2[0][2] = 1209ns;
slave_timing[0][9].t_rxd2[2][0] = 865ns;
slave_timing[0][9].t_rxd2[1][2] = 939ns;
slave_timing[0][9].t_rxd2[2][1] = 1206ns;

slave_timing[0][10].info_corner          = 1;
slave_timing[0][10].info_temp__j__       = 125;
slave_timing[0][10].info_i__quite_rec__  = 0.003000000;
slave_timing[0][10].info_dtr__ib__       = 1;
slave_timing[0][10].info_i__offset_rec__ = 0.000000000;
slave_timing[0][10].info_i__max_slave__  = 0.023000000;
slave_timing[0][10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][10].info_r__dsi_bus__    = 5.000;

slave_timing[0][10].t_rxd1[0][1] = 1100ns;
slave_timing[0][10].t_rxd1[1][0] = 1061ns;
slave_timing[0][10].t_rxd1[0][2] = 814ns;
slave_timing[0][10].t_rxd1[2][0] = 1310ns;
slave_timing[0][10].t_rxd2[0][2] = 1390ns;
slave_timing[0][10].t_rxd2[2][0] = 761ns;
slave_timing[0][10].t_rxd2[1][2] = 1166ns;
slave_timing[0][10].t_rxd2[2][1] = 981ns;

slave_timing[0][11].info_corner          = 1;
slave_timing[0][11].info_temp__j__       = 125;
slave_timing[0][11].info_i__quite_rec__  = 0.003000000;
slave_timing[0][11].info_dtr__ib__       = 1;
slave_timing[0][11].info_i__offset_rec__ = 0.000000000;
slave_timing[0][11].info_i__max_slave__  = 0.025000000;
slave_timing[0][11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][11].info_r__dsi_bus__    = 5.000;

slave_timing[0][11].t_rxd1[0][1] = 1053ns;
slave_timing[0][11].t_rxd1[1][0] = 1094ns;
slave_timing[0][11].t_rxd1[0][2] = 790ns;
slave_timing[0][11].t_rxd1[2][0] = 1335ns;
slave_timing[0][11].t_rxd2[0][2] = 1273ns;
slave_timing[0][11].t_rxd2[2][0] = 817ns;
slave_timing[0][11].t_rxd2[1][2] = 1030ns;
slave_timing[0][11].t_rxd2[2][1] = 1094ns;

slave_timing[0][12].info_corner          = 1;
slave_timing[0][12].info_temp__j__       = 125;
slave_timing[0][12].info_i__quite_rec__  = 0.003000000;
slave_timing[0][12].info_dtr__ib__       = -1;
slave_timing[0][12].info_i__offset_rec__ = 0.000000000;
slave_timing[0][12].info_i__max_slave__  = 0.023000000;
slave_timing[0][12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][12].info_r__dsi_bus__    = 5.000;

slave_timing[0][12].t_rxd1[0][1] = 1282ns;
slave_timing[0][12].t_rxd1[1][0] = 1254ns;
slave_timing[0][12].t_rxd1[0][2] = 953ns;
slave_timing[0][12].t_rxd1[2][0] = 1489ns;
slave_timing[0][12].t_rxd2[0][2] = 1360ns;
slave_timing[0][12].t_rxd2[2][0] = 855ns;
slave_timing[0][12].t_rxd2[1][2] = 1079ns;
slave_timing[0][12].t_rxd2[2][1] = 1098ns;

slave_timing[0][13].info_corner          = 1;
slave_timing[0][13].info_temp__j__       = 125;
slave_timing[0][13].info_i__quite_rec__  = 0.003000000;
slave_timing[0][13].info_dtr__ib__       = -1;
slave_timing[0][13].info_i__offset_rec__ = 0.000000000;
slave_timing[0][13].info_i__max_slave__  = 0.025000000;
slave_timing[0][13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][13].info_r__dsi_bus__    = 5.000;

slave_timing[0][13].t_rxd1[0][1] = 1226ns;
slave_timing[0][13].t_rxd1[1][0] = 1285ns;
slave_timing[0][13].t_rxd1[0][2] = 925ns;
slave_timing[0][13].t_rxd1[2][0] = 1514ns;
slave_timing[0][13].t_rxd2[0][2] = 1272ns;
slave_timing[0][13].t_rxd2[2][0] = 902ns;
slave_timing[0][13].t_rxd2[1][2] = 968ns;
slave_timing[0][13].t_rxd2[2][1] = 1228ns;

slave_timing[0][14].info_corner          = 1;
slave_timing[0][14].info_temp__j__       = 125;
slave_timing[0][14].info_i__quite_rec__  = 0.003000000;
slave_timing[0][14].info_dtr__ib__       = 1;
slave_timing[0][14].info_i__offset_rec__ = 0.000000000;
slave_timing[0][14].info_i__max_slave__  = 0.023000000;
slave_timing[0][14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][14].info_r__dsi_bus__    = 5.000;

slave_timing[0][14].t_rxd1[0][1] = 1317ns;
slave_timing[0][14].t_rxd1[1][0] = 1206ns;
slave_timing[0][14].t_rxd1[0][2] = 962ns;
slave_timing[0][14].t_rxd1[2][0] = 1444ns;
slave_timing[0][14].t_rxd2[0][2] = 1444ns;
slave_timing[0][14].t_rxd2[2][0] = 798ns;
slave_timing[0][14].t_rxd2[1][2] = 1187ns;
slave_timing[0][14].t_rxd2[2][1] = 1012ns;

slave_timing[0][15].info_corner          = 1;
slave_timing[0][15].info_temp__j__       = 125;
slave_timing[0][15].info_i__quite_rec__  = 0.003000000;
slave_timing[0][15].info_dtr__ib__       = 1;
slave_timing[0][15].info_i__offset_rec__ = 0.000000000;
slave_timing[0][15].info_i__max_slave__  = 0.025000000;
slave_timing[0][15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][15].info_r__dsi_bus__    = 5.000;

slave_timing[0][15].t_rxd1[0][1] = 1256ns;
slave_timing[0][15].t_rxd1[1][0] = 1237ns;
slave_timing[0][15].t_rxd1[0][2] = 935ns;
slave_timing[0][15].t_rxd1[2][0] = 1468ns;
slave_timing[0][15].t_rxd2[0][2] = 1330ns;
slave_timing[0][15].t_rxd2[2][0] = 852ns;
slave_timing[0][15].t_rxd2[1][2] = 1054ns;
slave_timing[0][15].t_rxd2[2][1] = 1117ns;

slave_timing[0][16].info_corner          = 1;
slave_timing[0][16].info_temp__j__       = 125;
slave_timing[0][16].info_i__quite_rec__  = 0.000000000;
slave_timing[0][16].info_dtr__ib__       = -1;
slave_timing[0][16].info_i__offset_rec__ = 0.000000000;
slave_timing[0][16].info_i__max_slave__  = 0.023000000;
slave_timing[0][16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][16].info_r__dsi_bus__    = 5.000;

slave_timing[0][16].t_rxd1[0][1] = 1059ns;
slave_timing[0][16].t_rxd1[1][0] = 1084ns;
slave_timing[0][16].t_rxd1[0][2] = 794ns;
slave_timing[0][16].t_rxd1[2][0] = 1324ns;
slave_timing[0][16].t_rxd2[0][2] = 1285ns;
slave_timing[0][16].t_rxd2[2][0] = 806ns;
slave_timing[0][16].t_rxd2[1][2] = 1050ns;
slave_timing[0][16].t_rxd2[2][1] = 1068ns;

slave_timing[0][17].info_corner          = 1;
slave_timing[0][17].info_temp__j__       = 125;
slave_timing[0][17].info_i__quite_rec__  = 0.000000000;
slave_timing[0][17].info_dtr__ib__       = -1;
slave_timing[0][17].info_i__offset_rec__ = 0.000000000;
slave_timing[0][17].info_i__max_slave__  = 0.025000000;
slave_timing[0][17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][17].info_r__dsi_bus__    = 5.000;

slave_timing[0][17].t_rxd1[0][1] = 1017ns;
slave_timing[0][17].t_rxd1[1][0] = 1111ns;
slave_timing[0][17].t_rxd1[0][2] = 770ns;
slave_timing[0][17].t_rxd1[2][0] = 1348ns;
slave_timing[0][17].t_rxd2[0][2] = 1195ns;
slave_timing[0][17].t_rxd2[2][0] = 851ns;
slave_timing[0][17].t_rxd2[1][2] = 938ns;
slave_timing[0][17].t_rxd2[2][1] = 1187ns;

slave_timing[0][18].info_corner          = 1;
slave_timing[0][18].info_temp__j__       = 125;
slave_timing[0][18].info_i__quite_rec__  = 0.000000000;
slave_timing[0][18].info_dtr__ib__       = 1;
slave_timing[0][18].info_i__offset_rec__ = 0.000000000;
slave_timing[0][18].info_i__max_slave__  = 0.023000000;
slave_timing[0][18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][18].info_r__dsi_bus__    = 5.000;

slave_timing[0][18].t_rxd1[0][1] = 1097ns;
slave_timing[0][18].t_rxd1[1][0] = 1026ns;
slave_timing[0][18].t_rxd1[0][2] = 808ns;
slave_timing[0][18].t_rxd1[2][0] = 1266ns;
slave_timing[0][18].t_rxd2[0][2] = 1386ns;
slave_timing[0][18].t_rxd2[2][0] = 737ns;
slave_timing[0][18].t_rxd2[1][2] = 1178ns;
slave_timing[0][18].t_rxd2[2][1] = 941ns;

slave_timing[0][19].info_corner          = 1;
slave_timing[0][19].info_temp__j__       = 125;
slave_timing[0][19].info_i__quite_rec__  = 0.000000000;
slave_timing[0][19].info_dtr__ib__       = 1;
slave_timing[0][19].info_i__offset_rec__ = 0.000000000;
slave_timing[0][19].info_i__max_slave__  = 0.025000000;
slave_timing[0][19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][19].info_r__dsi_bus__    = 5.000;

slave_timing[0][19].t_rxd1[0][1] = 1048ns;
slave_timing[0][19].t_rxd1[1][0] = 1058ns;
slave_timing[0][19].t_rxd1[0][2] = 775ns;
slave_timing[0][19].t_rxd1[2][0] = 1292ns;
slave_timing[0][19].t_rxd2[0][2] = 1248ns;
slave_timing[0][19].t_rxd2[2][0] = 794ns;
slave_timing[0][19].t_rxd2[1][2] = 1038ns;
slave_timing[0][19].t_rxd2[2][1] = 1051ns;

slave_timing[0][20].info_corner          = 1;
slave_timing[0][20].info_temp__j__       = 125;
slave_timing[0][20].info_i__quite_rec__  = 0.000000000;
slave_timing[0][20].info_dtr__ib__       = -1;
slave_timing[0][20].info_i__offset_rec__ = 0.000000000;
slave_timing[0][20].info_i__max_slave__  = 0.023000000;
slave_timing[0][20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][20].info_r__dsi_bus__    = 5.000;

slave_timing[0][20].t_rxd1[0][1] = 1283ns;
slave_timing[0][20].t_rxd1[1][0] = 1227ns;
slave_timing[0][20].t_rxd1[0][2] = 954ns;
slave_timing[0][20].t_rxd1[2][0] = 1455ns;
slave_timing[0][20].t_rxd2[0][2] = 1340ns;
slave_timing[0][20].t_rxd2[2][0] = 843ns;
slave_timing[0][20].t_rxd2[1][2] = 1073ns;
slave_timing[0][20].t_rxd2[2][1] = 1093ns;

slave_timing[0][21].info_corner          = 1;
slave_timing[0][21].info_temp__j__       = 125;
slave_timing[0][21].info_i__quite_rec__  = 0.000000000;
slave_timing[0][21].info_dtr__ib__       = -1;
slave_timing[0][21].info_i__offset_rec__ = 0.000000000;
slave_timing[0][21].info_i__max_slave__  = 0.025000000;
slave_timing[0][21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][21].info_r__dsi_bus__    = 5.000;

slave_timing[0][21].t_rxd1[0][1] = 1227ns;
slave_timing[0][21].t_rxd1[1][0] = 1256ns;
slave_timing[0][21].t_rxd1[0][2] = 928ns;
slave_timing[0][21].t_rxd1[2][0] = 1480ns;
slave_timing[0][21].t_rxd2[0][2] = 1257ns;
slave_timing[0][21].t_rxd2[2][0] = 890ns;
slave_timing[0][21].t_rxd2[1][2] = 964ns;
slave_timing[0][21].t_rxd2[2][1] = 1203ns;

slave_timing[0][22].info_corner          = 1;
slave_timing[0][22].info_temp__j__       = 125;
slave_timing[0][22].info_i__quite_rec__  = 0.000000000;
slave_timing[0][22].info_dtr__ib__       = 1;
slave_timing[0][22].info_i__offset_rec__ = 0.000000000;
slave_timing[0][22].info_i__max_slave__  = 0.023000000;
slave_timing[0][22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][22].info_r__dsi_bus__    = 5.000;

slave_timing[0][22].t_rxd1[0][1] = 1339ns;
slave_timing[0][22].t_rxd1[1][0] = 1168ns;
slave_timing[0][22].t_rxd1[0][2] = 974ns;
slave_timing[0][22].t_rxd1[2][0] = 1397ns;
slave_timing[0][22].t_rxd2[0][2] = 1439ns;
slave_timing[0][22].t_rxd2[2][0] = 772ns;
slave_timing[0][22].t_rxd2[1][2] = 1195ns;
slave_timing[0][22].t_rxd2[2][1] = 969ns;

slave_timing[0][23].info_corner          = 1;
slave_timing[0][23].info_temp__j__       = 125;
slave_timing[0][23].info_i__quite_rec__  = 0.000000000;
slave_timing[0][23].info_dtr__ib__       = 1;
slave_timing[0][23].info_i__offset_rec__ = 0.000000000;
slave_timing[0][23].info_i__max_slave__  = 0.025000000;
slave_timing[0][23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][23].info_r__dsi_bus__    = 5.000;

slave_timing[0][23].t_rxd1[0][1] = 1278ns;
slave_timing[0][23].t_rxd1[1][0] = 1199ns;
slave_timing[0][23].t_rxd1[0][2] = 946ns;
slave_timing[0][23].t_rxd1[2][0] = 1424ns;
slave_timing[0][23].t_rxd2[0][2] = 1320ns;
slave_timing[0][23].t_rxd2[2][0] = 830ns;
slave_timing[0][23].t_rxd2[1][2] = 1058ns;
slave_timing[0][23].t_rxd2[2][1] = 1076ns;

slave_timing[0][24].info_corner          = 1;
slave_timing[0][24].info_temp__j__       = 125;
slave_timing[0][24].info_i__quite_rec__  = 0.040000000;
slave_timing[0][24].info_dtr__ib__       = -1;
slave_timing[0][24].info_i__offset_rec__ = 0.000000000;
slave_timing[0][24].info_i__max_slave__  = 0.023000000;
slave_timing[0][24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][24].info_r__dsi_bus__    = 5.000;

slave_timing[0][24].t_rxd1[0][1] = 1094ns;
slave_timing[0][24].t_rxd1[1][0] = 1110ns;
slave_timing[0][24].t_rxd1[0][2] = 807ns;
slave_timing[0][24].t_rxd1[2][0] = 1371ns;
slave_timing[0][24].t_rxd2[0][2] = 1312ns;
slave_timing[0][24].t_rxd2[2][0] = 821ns;
slave_timing[0][24].t_rxd2[1][2] = 1074ns;
slave_timing[0][24].t_rxd2[2][1] = 1082ns;

slave_timing[0][25].info_corner          = 1;
slave_timing[0][25].info_temp__j__       = 125;
slave_timing[0][25].info_i__quite_rec__  = 0.040000000;
slave_timing[0][25].info_dtr__ib__       = -1;
slave_timing[0][25].info_i__offset_rec__ = 0.000000000;
slave_timing[0][25].info_i__max_slave__  = 0.025000000;
slave_timing[0][25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][25].info_r__dsi_bus__    = 5.000;

slave_timing[0][25].t_rxd1[0][1] = 1034ns;
slave_timing[0][25].t_rxd1[1][0] = 1154ns;
slave_timing[0][25].t_rxd1[0][2] = 785ns;
slave_timing[0][25].t_rxd1[2][0] = 1401ns;
slave_timing[0][25].t_rxd2[0][2] = 1224ns;
slave_timing[0][25].t_rxd2[2][0] = 871ns;
slave_timing[0][25].t_rxd2[1][2] = 943ns;
slave_timing[0][25].t_rxd2[2][1] = 1224ns;

slave_timing[0][26].info_corner          = 1;
slave_timing[0][26].info_temp__j__       = 125;
slave_timing[0][26].info_i__quite_rec__  = 0.040000000;
slave_timing[0][26].info_dtr__ib__       = 1;
slave_timing[0][26].info_i__offset_rec__ = 0.000000000;
slave_timing[0][26].info_i__max_slave__  = 0.023000000;
slave_timing[0][26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][26].info_r__dsi_bus__    = 5.000;

slave_timing[0][26].t_rxd1[0][1] = 1125ns;
slave_timing[0][26].t_rxd1[1][0] = 1075ns;
slave_timing[0][26].t_rxd1[0][2] = 828ns;
slave_timing[0][26].t_rxd1[2][0] = 1333ns;
slave_timing[0][26].t_rxd2[0][2] = 1420ns;
slave_timing[0][26].t_rxd2[2][0] = 768ns;
slave_timing[0][26].t_rxd2[1][2] = 1180ns;
slave_timing[0][26].t_rxd2[2][1] = 994ns;

slave_timing[0][27].info_corner          = 1;
slave_timing[0][27].info_temp__j__       = 125;
slave_timing[0][27].info_i__quite_rec__  = 0.040000000;
slave_timing[0][27].info_dtr__ib__       = 1;
slave_timing[0][27].info_i__offset_rec__ = 0.000000000;
slave_timing[0][27].info_i__max_slave__  = 0.025000000;
slave_timing[0][27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][27].info_r__dsi_bus__    = 5.000;

slave_timing[0][27].t_rxd1[0][1] = 1075ns;
slave_timing[0][27].t_rxd1[1][0] = 1108ns;
slave_timing[0][27].t_rxd1[0][2] = 803ns;
slave_timing[0][27].t_rxd1[2][0] = 1362ns;
slave_timing[0][27].t_rxd2[0][2] = 1300ns;
slave_timing[0][27].t_rxd2[2][0] = 824ns;
slave_timing[0][27].t_rxd2[1][2] = 1045ns;
slave_timing[0][27].t_rxd2[2][1] = 1109ns;

slave_timing[0][28].info_corner          = 1;
slave_timing[0][28].info_temp__j__       = 125;
slave_timing[0][28].info_i__quite_rec__  = 0.040000000;
slave_timing[0][28].info_dtr__ib__       = -1;
slave_timing[0][28].info_i__offset_rec__ = 0.000000000;
slave_timing[0][28].info_i__max_slave__  = 0.023000000;
slave_timing[0][28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][28].info_r__dsi_bus__    = 5.000;

slave_timing[0][28].t_rxd1[0][1] = 1191ns;
slave_timing[0][28].t_rxd1[1][0] = 1225ns;
slave_timing[0][28].t_rxd1[0][2] = 904ns;
slave_timing[0][28].t_rxd1[2][0] = 1459ns;
slave_timing[0][28].t_rxd2[0][2] = 1362ns;
slave_timing[0][28].t_rxd2[2][0] = 868ns;
slave_timing[0][28].t_rxd2[1][2] = 1104ns;
slave_timing[0][28].t_rxd2[2][1] = 1125ns;

slave_timing[0][29].info_corner          = 1;
slave_timing[0][29].info_temp__j__       = 125;
slave_timing[0][29].info_i__quite_rec__  = 0.040000000;
slave_timing[0][29].info_dtr__ib__       = -1;
slave_timing[0][29].info_i__offset_rec__ = 0.000000000;
slave_timing[0][29].info_i__max_slave__  = 0.025000000;
slave_timing[0][29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][29].info_r__dsi_bus__    = 5.000;

slave_timing[0][29].t_rxd1[0][1] = 1143ns;
slave_timing[0][29].t_rxd1[1][0] = 1254ns;
slave_timing[0][29].t_rxd1[0][2] = 879ns;
slave_timing[0][29].t_rxd1[2][0] = 1483ns;
slave_timing[0][29].t_rxd2[0][2] = 1284ns;
slave_timing[0][29].t_rxd2[2][0] = 912ns;
slave_timing[0][29].t_rxd2[1][2] = 994ns;
slave_timing[0][29].t_rxd2[2][1] = 1214ns;

slave_timing[0][30].info_corner          = 1;
slave_timing[0][30].info_temp__j__       = 125;
slave_timing[0][30].info_i__quite_rec__  = 0.040000000;
slave_timing[0][30].info_dtr__ib__       = 1;
slave_timing[0][30].info_i__offset_rec__ = 0.000000000;
slave_timing[0][30].info_i__max_slave__  = 0.023000000;
slave_timing[0][30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][30].info_r__dsi_bus__    = 5.000;

slave_timing[0][30].t_rxd1[0][1] = 1236ns;
slave_timing[0][30].t_rxd1[1][0] = 1170ns;
slave_timing[0][30].t_rxd1[0][2] = 922ns;
slave_timing[0][30].t_rxd1[2][0] = 1415ns;
slave_timing[0][30].t_rxd2[0][2] = 1453ns;
slave_timing[0][30].t_rxd2[2][0] = 814ns;
slave_timing[0][30].t_rxd2[1][2] = 1219ns;
slave_timing[0][30].t_rxd2[2][1] = 1029ns;

slave_timing[0][31].info_corner          = 1;
slave_timing[0][31].info_temp__j__       = 125;
slave_timing[0][31].info_i__quite_rec__  = 0.040000000;
slave_timing[0][31].info_dtr__ib__       = 1;
slave_timing[0][31].info_i__offset_rec__ = 0.000000000;
slave_timing[0][31].info_i__max_slave__  = 0.025000000;
slave_timing[0][31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][31].info_r__dsi_bus__    = 5.000;

slave_timing[0][31].t_rxd1[0][1] = 1183ns;
slave_timing[0][31].t_rxd1[1][0] = 1204ns;
slave_timing[0][31].t_rxd1[0][2] = 896ns;
slave_timing[0][31].t_rxd1[2][0] = 1442ns;
slave_timing[0][31].t_rxd2[0][2] = 1350ns;
slave_timing[0][31].t_rxd2[2][0] = 867ns;
slave_timing[0][31].t_rxd2[1][2] = 1089ns;
slave_timing[0][31].t_rxd2[2][1] = 1130ns;


slave_timing[1][192+0].info_corner          = 3;
slave_timing[1][192+0].info_temp__j__       = -40;
slave_timing[1][192+0].info_i__quite_rec__  = 0.006000000;
slave_timing[1][192+0].info_dtr__ib__       = -1;
slave_timing[1][192+0].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+0].info_i__max_slave__  = 0.023000000;
slave_timing[1][192+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][192+0].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+0].t_rxd1[0][1] = 1653ns;
slave_timing[1][192+0].t_rxd1[1][0] = 1671ns;
slave_timing[1][192+0].t_rxd1[0][2] = 1243ns;
slave_timing[1][192+0].t_rxd1[2][0] = 2030ns;
slave_timing[1][192+0].t_rxd2[0][2] = 1992ns;
slave_timing[1][192+0].t_rxd2[2][0] = 1258ns;
slave_timing[1][192+0].t_rxd2[1][2] = 1624ns;
slave_timing[1][192+0].t_rxd2[2][1] = 1666ns;

slave_timing[1][192+1].info_corner          = 3;
slave_timing[1][192+1].info_temp__j__       = -40;
slave_timing[1][192+1].info_i__quite_rec__  = 0.006000000;
slave_timing[1][192+1].info_dtr__ib__       = -1;
slave_timing[1][192+1].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+1].info_i__max_slave__  = 0.025000000;
slave_timing[1][192+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][192+1].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+1].t_rxd1[0][1] = 1591ns;
slave_timing[1][192+1].t_rxd1[1][0] = 1718ns;
slave_timing[1][192+1].t_rxd1[0][2] = 1212ns;
slave_timing[1][192+1].t_rxd1[2][0] = 2065ns;
slave_timing[1][192+1].t_rxd2[0][2] = 1877ns;
slave_timing[1][192+1].t_rxd2[2][0] = 1338ns;
slave_timing[1][192+1].t_rxd2[1][2] = 1453ns;
slave_timing[1][192+1].t_rxd2[2][1] = 1845ns;

slave_timing[1][192+2].info_corner          = 3;
slave_timing[1][192+2].info_temp__j__       = -40;
slave_timing[1][192+2].info_i__quite_rec__  = 0.006000000;
slave_timing[1][192+2].info_dtr__ib__       = 1;
slave_timing[1][192+2].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+2].info_i__max_slave__  = 0.023000000;
slave_timing[1][192+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][192+2].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+2].t_rxd1[0][1] = 1703ns;
slave_timing[1][192+2].t_rxd1[1][0] = 1631ns;
slave_timing[1][192+2].t_rxd1[0][2] = 1270ns;
slave_timing[1][192+2].t_rxd1[2][0] = 2002ns;
slave_timing[1][192+2].t_rxd2[0][2] = 2099ns;
slave_timing[1][192+2].t_rxd2[2][0] = 1184ns;
slave_timing[1][192+2].t_rxd2[1][2] = 1771ns;
slave_timing[1][192+2].t_rxd2[2][1] = 1540ns;

slave_timing[1][192+3].info_corner          = 3;
slave_timing[1][192+3].info_temp__j__       = -40;
slave_timing[1][192+3].info_i__quite_rec__  = 0.006000000;
slave_timing[1][192+3].info_dtr__ib__       = 1;
slave_timing[1][192+3].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+3].info_i__max_slave__  = 0.025000000;
slave_timing[1][192+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][192+3].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+3].t_rxd1[0][1] = 1634ns;
slave_timing[1][192+3].t_rxd1[1][0] = 1682ns;
slave_timing[1][192+3].t_rxd1[0][2] = 1233ns;
slave_timing[1][192+3].t_rxd1[2][0] = 2038ns;
slave_timing[1][192+3].t_rxd2[0][2] = 1957ns;
slave_timing[1][192+3].t_rxd2[2][0] = 1274ns;
slave_timing[1][192+3].t_rxd2[1][2] = 1577ns;
slave_timing[1][192+3].t_rxd2[2][1] = 1712ns;

slave_timing[1][192+4].info_corner          = 3;
slave_timing[1][192+4].info_temp__j__       = -40;
slave_timing[1][192+4].info_i__quite_rec__  = 0.006000000;
slave_timing[1][192+4].info_dtr__ib__       = -1;
slave_timing[1][192+4].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+4].info_i__max_slave__  = 0.023000000;
slave_timing[1][192+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][192+4].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+4].t_rxd1[0][1] = 1737ns;
slave_timing[1][192+4].t_rxd1[1][0] = 1747ns;
slave_timing[1][192+4].t_rxd1[0][2] = 1313ns;
slave_timing[1][192+4].t_rxd1[2][0] = 2103ns;
slave_timing[1][192+4].t_rxd2[0][2] = 2013ns;
slave_timing[1][192+4].t_rxd2[2][0] = 1275ns;
slave_timing[1][192+4].t_rxd2[1][2] = 1638ns;
slave_timing[1][192+4].t_rxd2[2][1] = 1685ns;

slave_timing[1][192+5].info_corner          = 3;
slave_timing[1][192+5].info_temp__j__       = -40;
slave_timing[1][192+5].info_i__quite_rec__  = 0.006000000;
slave_timing[1][192+5].info_dtr__ib__       = -1;
slave_timing[1][192+5].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+5].info_i__max_slave__  = 0.025000000;
slave_timing[1][192+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][192+5].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+5].t_rxd1[0][1] = 1671ns;
slave_timing[1][192+5].t_rxd1[1][0] = 1796ns;
slave_timing[1][192+5].t_rxd1[0][2] = 1278ns;
slave_timing[1][192+5].t_rxd1[2][0] = 2136ns;
slave_timing[1][192+5].t_rxd2[0][2] = 1897ns;
slave_timing[1][192+5].t_rxd2[2][0] = 1356ns;
slave_timing[1][192+5].t_rxd2[1][2] = 1465ns;
slave_timing[1][192+5].t_rxd2[2][1] = 1857ns;

slave_timing[1][192+6].info_corner          = 3;
slave_timing[1][192+6].info_temp__j__       = -40;
slave_timing[1][192+6].info_i__quite_rec__  = 0.006000000;
slave_timing[1][192+6].info_dtr__ib__       = 1;
slave_timing[1][192+6].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+6].info_i__max_slave__  = 0.023000000;
slave_timing[1][192+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][192+6].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+6].t_rxd1[0][1] = 1776ns;
slave_timing[1][192+6].t_rxd1[1][0] = 1703ns;
slave_timing[1][192+6].t_rxd1[0][2] = 1333ns;
slave_timing[1][192+6].t_rxd1[2][0] = 2071ns;
slave_timing[1][192+6].t_rxd2[0][2] = 2118ns;
slave_timing[1][192+6].t_rxd2[2][0] = 1202ns;
slave_timing[1][192+6].t_rxd2[1][2] = 1783ns;
slave_timing[1][192+6].t_rxd2[2][1] = 1554ns;

slave_timing[1][192+7].info_corner          = 3;
slave_timing[1][192+7].info_temp__j__       = -40;
slave_timing[1][192+7].info_i__quite_rec__  = 0.006000000;
slave_timing[1][192+7].info_dtr__ib__       = 1;
slave_timing[1][192+7].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+7].info_i__max_slave__  = 0.025000000;
slave_timing[1][192+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][192+7].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+7].t_rxd1[0][1] = 1708ns;
slave_timing[1][192+7].t_rxd1[1][0] = 1751ns;
slave_timing[1][192+7].t_rxd1[0][2] = 1294ns;
slave_timing[1][192+7].t_rxd1[2][0] = 2105ns;
slave_timing[1][192+7].t_rxd2[0][2] = 1977ns;
slave_timing[1][192+7].t_rxd2[2][0] = 1293ns;
slave_timing[1][192+7].t_rxd2[1][2] = 1589ns;
slave_timing[1][192+7].t_rxd2[2][1] = 1725ns;

slave_timing[1][192+8].info_corner          = 3;
slave_timing[1][192+8].info_temp__j__       = -40;
slave_timing[1][192+8].info_i__quite_rec__  = 0.003000000;
slave_timing[1][192+8].info_dtr__ib__       = -1;
slave_timing[1][192+8].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+8].info_i__max_slave__  = 0.023000000;
slave_timing[1][192+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][192+8].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+8].t_rxd1[0][1] = 1648ns;
slave_timing[1][192+8].t_rxd1[1][0] = 1682ns;
slave_timing[1][192+8].t_rxd1[0][2] = 1241ns;
slave_timing[1][192+8].t_rxd1[2][0] = 2039ns;
slave_timing[1][192+8].t_rxd2[0][2] = 1985ns;
slave_timing[1][192+8].t_rxd2[2][0] = 1257ns;
slave_timing[1][192+8].t_rxd2[1][2] = 1615ns;
slave_timing[1][192+8].t_rxd2[2][1] = 1675ns;

slave_timing[1][192+9].info_corner          = 3;
slave_timing[1][192+9].info_temp__j__       = -40;
slave_timing[1][192+9].info_i__quite_rec__  = 0.003000000;
slave_timing[1][192+9].info_dtr__ib__       = -1;
slave_timing[1][192+9].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+9].info_i__max_slave__  = 0.025000000;
slave_timing[1][192+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][192+9].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+9].t_rxd1[0][1] = 1586ns;
slave_timing[1][192+9].t_rxd1[1][0] = 1730ns;
slave_timing[1][192+9].t_rxd1[0][2] = 1209ns;
slave_timing[1][192+9].t_rxd1[2][0] = 2075ns;
slave_timing[1][192+9].t_rxd2[0][2] = 1870ns;
slave_timing[1][192+9].t_rxd2[2][0] = 1339ns;
slave_timing[1][192+9].t_rxd2[1][2] = 1444ns;
slave_timing[1][192+9].t_rxd2[2][1] = 1849ns;

slave_timing[1][192+10].info_corner          = 3;
slave_timing[1][192+10].info_temp__j__       = -40;
slave_timing[1][192+10].info_i__quite_rec__  = 0.003000000;
slave_timing[1][192+10].info_dtr__ib__       = 1;
slave_timing[1][192+10].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+10].info_i__max_slave__  = 0.023000000;
slave_timing[1][192+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][192+10].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+10].t_rxd1[0][1] = 1695ns;
slave_timing[1][192+10].t_rxd1[1][0] = 1638ns;
slave_timing[1][192+10].t_rxd1[0][2] = 1266ns;
slave_timing[1][192+10].t_rxd1[2][0] = 2006ns;
slave_timing[1][192+10].t_rxd2[0][2] = 2093ns;
slave_timing[1][192+10].t_rxd2[2][0] = 1190ns;
slave_timing[1][192+10].t_rxd2[1][2] = 1764ns;
slave_timing[1][192+10].t_rxd2[2][1] = 1549ns;

slave_timing[1][192+11].info_corner          = 3;
slave_timing[1][192+11].info_temp__j__       = -40;
slave_timing[1][192+11].info_i__quite_rec__  = 0.003000000;
slave_timing[1][192+11].info_dtr__ib__       = 1;
slave_timing[1][192+11].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+11].info_i__max_slave__  = 0.025000000;
slave_timing[1][192+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][192+11].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+11].t_rxd1[0][1] = 1626ns;
slave_timing[1][192+11].t_rxd1[1][0] = 1685ns;
slave_timing[1][192+11].t_rxd1[0][2] = 1229ns;
slave_timing[1][192+11].t_rxd1[2][0] = 2040ns;
slave_timing[1][192+11].t_rxd2[0][2] = 1953ns;
slave_timing[1][192+11].t_rxd2[2][0] = 1278ns;
slave_timing[1][192+11].t_rxd2[1][2] = 1569ns;
slave_timing[1][192+11].t_rxd2[2][1] = 1720ns;

slave_timing[1][192+12].info_corner          = 3;
slave_timing[1][192+12].info_temp__j__       = -40;
slave_timing[1][192+12].info_i__quite_rec__  = 0.003000000;
slave_timing[1][192+12].info_dtr__ib__       = -1;
slave_timing[1][192+12].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+12].info_i__max_slave__  = 0.023000000;
slave_timing[1][192+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][192+12].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+12].t_rxd1[0][1] = 1731ns;
slave_timing[1][192+12].t_rxd1[1][0] = 1761ns;
slave_timing[1][192+12].t_rxd1[0][2] = 1313ns;
slave_timing[1][192+12].t_rxd1[2][0] = 2114ns;
slave_timing[1][192+12].t_rxd2[0][2] = 2007ns;
slave_timing[1][192+12].t_rxd2[2][0] = 1277ns;
slave_timing[1][192+12].t_rxd2[1][2] = 1653ns;
slave_timing[1][192+12].t_rxd2[2][1] = 1664ns;

slave_timing[1][192+13].info_corner          = 3;
slave_timing[1][192+13].info_temp__j__       = -40;
slave_timing[1][192+13].info_i__quite_rec__  = 0.003000000;
slave_timing[1][192+13].info_dtr__ib__       = -1;
slave_timing[1][192+13].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+13].info_i__max_slave__  = 0.025000000;
slave_timing[1][192+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][192+13].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+13].t_rxd1[0][1] = 1667ns;
slave_timing[1][192+13].t_rxd1[1][0] = 1807ns;
slave_timing[1][192+13].t_rxd1[0][2] = 1276ns;
slave_timing[1][192+13].t_rxd1[2][0] = 2148ns;
slave_timing[1][192+13].t_rxd2[0][2] = 1892ns;
slave_timing[1][192+13].t_rxd2[2][0] = 1357ns;
slave_timing[1][192+13].t_rxd2[1][2] = 1458ns;
slave_timing[1][192+13].t_rxd2[2][1] = 1859ns;

slave_timing[1][192+14].info_corner          = 3;
slave_timing[1][192+14].info_temp__j__       = -40;
slave_timing[1][192+14].info_i__quite_rec__  = 0.003000000;
slave_timing[1][192+14].info_dtr__ib__       = 1;
slave_timing[1][192+14].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+14].info_i__max_slave__  = 0.023000000;
slave_timing[1][192+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][192+14].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+14].t_rxd1[0][1] = 1773ns;
slave_timing[1][192+14].t_rxd1[1][0] = 1707ns;
slave_timing[1][192+14].t_rxd1[0][2] = 1330ns;
slave_timing[1][192+14].t_rxd1[2][0] = 2073ns;
slave_timing[1][192+14].t_rxd2[0][2] = 2110ns;
slave_timing[1][192+14].t_rxd2[2][0] = 1200ns;
slave_timing[1][192+14].t_rxd2[1][2] = 1773ns;
slave_timing[1][192+14].t_rxd2[2][1] = 1559ns;

slave_timing[1][192+15].info_corner          = 3;
slave_timing[1][192+15].info_temp__j__       = -40;
slave_timing[1][192+15].info_i__quite_rec__  = 0.003000000;
slave_timing[1][192+15].info_dtr__ib__       = 1;
slave_timing[1][192+15].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+15].info_i__max_slave__  = 0.025000000;
slave_timing[1][192+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][192+15].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+15].t_rxd1[0][1] = 1703ns;
slave_timing[1][192+15].t_rxd1[1][0] = 1759ns;
slave_timing[1][192+15].t_rxd1[0][2] = 1293ns;
slave_timing[1][192+15].t_rxd1[2][0] = 2109ns;
slave_timing[1][192+15].t_rxd2[0][2] = 1972ns;
slave_timing[1][192+15].t_rxd2[2][0] = 1294ns;
slave_timing[1][192+15].t_rxd2[1][2] = 1582ns;
slave_timing[1][192+15].t_rxd2[2][1] = 1727ns;

slave_timing[1][192+16].info_corner          = 3;
slave_timing[1][192+16].info_temp__j__       = -40;
slave_timing[1][192+16].info_i__quite_rec__  = 0.000000000;
slave_timing[1][192+16].info_dtr__ib__       = -1;
slave_timing[1][192+16].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+16].info_i__max_slave__  = 0.023000000;
slave_timing[1][192+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][192+16].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+16].t_rxd1[0][1] = 1664ns;
slave_timing[1][192+16].t_rxd1[1][0] = 1663ns;
slave_timing[1][192+16].t_rxd1[0][2] = 1253ns;
slave_timing[1][192+16].t_rxd1[2][0] = 2024ns;
slave_timing[1][192+16].t_rxd2[0][2] = 1999ns;
slave_timing[1][192+16].t_rxd2[2][0] = 1251ns;
slave_timing[1][192+16].t_rxd2[1][2] = 1631ns;
slave_timing[1][192+16].t_rxd2[2][1] = 1660ns;

slave_timing[1][192+17].info_corner          = 3;
slave_timing[1][192+17].info_temp__j__       = -40;
slave_timing[1][192+17].info_i__quite_rec__  = 0.000000000;
slave_timing[1][192+17].info_dtr__ib__       = -1;
slave_timing[1][192+17].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+17].info_i__max_slave__  = 0.025000000;
slave_timing[1][192+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][192+17].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+17].t_rxd1[0][1] = 1600ns;
slave_timing[1][192+17].t_rxd1[1][0] = 1709ns;
slave_timing[1][192+17].t_rxd1[0][2] = 1216ns;
slave_timing[1][192+17].t_rxd1[2][0] = 2059ns;
slave_timing[1][192+17].t_rxd2[0][2] = 1879ns;
slave_timing[1][192+17].t_rxd2[2][0] = 1332ns;
slave_timing[1][192+17].t_rxd2[1][2] = 1456ns;
slave_timing[1][192+17].t_rxd2[2][1] = 1833ns;

slave_timing[1][192+18].info_corner          = 3;
slave_timing[1][192+18].info_temp__j__       = -40;
slave_timing[1][192+18].info_i__quite_rec__  = 0.000000000;
slave_timing[1][192+18].info_dtr__ib__       = 1;
slave_timing[1][192+18].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+18].info_i__max_slave__  = 0.023000000;
slave_timing[1][192+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][192+18].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+18].t_rxd1[0][1] = 1714ns;
slave_timing[1][192+18].t_rxd1[1][0] = 1618ns;
slave_timing[1][192+18].t_rxd1[0][2] = 1276ns;
slave_timing[1][192+18].t_rxd1[2][0] = 1994ns;
slave_timing[1][192+18].t_rxd2[0][2] = 2107ns;
slave_timing[1][192+18].t_rxd2[2][0] = 1177ns;
slave_timing[1][192+18].t_rxd2[1][2] = 1781ns;
slave_timing[1][192+18].t_rxd2[2][1] = 1526ns;

slave_timing[1][192+19].info_corner          = 3;
slave_timing[1][192+19].info_temp__j__       = -40;
slave_timing[1][192+19].info_i__quite_rec__  = 0.000000000;
slave_timing[1][192+19].info_dtr__ib__       = 1;
slave_timing[1][192+19].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+19].info_i__max_slave__  = 0.025000000;
slave_timing[1][192+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][192+19].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+19].t_rxd1[0][1] = 1645ns;
slave_timing[1][192+19].t_rxd1[1][0] = 1672ns;
slave_timing[1][192+19].t_rxd1[0][2] = 1239ns;
slave_timing[1][192+19].t_rxd1[2][0] = 2031ns;
slave_timing[1][192+19].t_rxd2[0][2] = 1964ns;
slave_timing[1][192+19].t_rxd2[2][0] = 1270ns;
slave_timing[1][192+19].t_rxd2[1][2] = 1587ns;
slave_timing[1][192+19].t_rxd2[2][1] = 1698ns;

slave_timing[1][192+20].info_corner          = 3;
slave_timing[1][192+20].info_temp__j__       = -40;
slave_timing[1][192+20].info_i__quite_rec__  = 0.000000000;
slave_timing[1][192+20].info_dtr__ib__       = -1;
slave_timing[1][192+20].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+20].info_i__max_slave__  = 0.023000000;
slave_timing[1][192+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][192+20].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+20].t_rxd1[0][1] = 1750ns;
slave_timing[1][192+20].t_rxd1[1][0] = 1738ns;
slave_timing[1][192+20].t_rxd1[0][2] = 1323ns;
slave_timing[1][192+20].t_rxd1[2][0] = 2098ns;
slave_timing[1][192+20].t_rxd2[0][2] = 2018ns;
slave_timing[1][192+20].t_rxd2[2][0] = 1266ns;
slave_timing[1][192+20].t_rxd2[1][2] = 1645ns;
slave_timing[1][192+20].t_rxd2[2][1] = 1644ns;

slave_timing[1][192+21].info_corner          = 3;
slave_timing[1][192+21].info_temp__j__       = -40;
slave_timing[1][192+21].info_i__quite_rec__  = 0.000000000;
slave_timing[1][192+21].info_dtr__ib__       = -1;
slave_timing[1][192+21].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+21].info_i__max_slave__  = 0.025000000;
slave_timing[1][192+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][192+21].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+21].t_rxd1[0][1] = 1685ns;
slave_timing[1][192+21].t_rxd1[1][0] = 1785ns;
slave_timing[1][192+21].t_rxd1[0][2] = 1287ns;
slave_timing[1][192+21].t_rxd1[2][0] = 2133ns;
slave_timing[1][192+21].t_rxd2[0][2] = 1901ns;
slave_timing[1][192+21].t_rxd2[2][0] = 1350ns;
slave_timing[1][192+21].t_rxd2[1][2] = 1470ns;
slave_timing[1][192+21].t_rxd2[2][1] = 1844ns;

slave_timing[1][192+22].info_corner          = 3;
slave_timing[1][192+22].info_temp__j__       = -40;
slave_timing[1][192+22].info_i__quite_rec__  = 0.000000000;
slave_timing[1][192+22].info_dtr__ib__       = 1;
slave_timing[1][192+22].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+22].info_i__max_slave__  = 0.023000000;
slave_timing[1][192+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][192+22].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+22].t_rxd1[0][1] = 1795ns;
slave_timing[1][192+22].t_rxd1[1][0] = 1691ns;
slave_timing[1][192+22].t_rxd1[0][2] = 1342ns;
slave_timing[1][192+22].t_rxd1[2][0] = 2063ns;
slave_timing[1][192+22].t_rxd2[0][2] = 2124ns;
slave_timing[1][192+22].t_rxd2[2][0] = 1191ns;
slave_timing[1][192+22].t_rxd2[1][2] = 1793ns;
slave_timing[1][192+22].t_rxd2[2][1] = 1540ns;

slave_timing[1][192+23].info_corner          = 3;
slave_timing[1][192+23].info_temp__j__       = -40;
slave_timing[1][192+23].info_i__quite_rec__  = 0.000000000;
slave_timing[1][192+23].info_dtr__ib__       = 1;
slave_timing[1][192+23].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+23].info_i__max_slave__  = 0.025000000;
slave_timing[1][192+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][192+23].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+23].t_rxd1[0][1] = 1724ns;
slave_timing[1][192+23].t_rxd1[1][0] = 1741ns;
slave_timing[1][192+23].t_rxd1[0][2] = 1304ns;
slave_timing[1][192+23].t_rxd1[2][0] = 2098ns;
slave_timing[1][192+23].t_rxd2[0][2] = 1982ns;
slave_timing[1][192+23].t_rxd2[2][0] = 1286ns;
slave_timing[1][192+23].t_rxd2[1][2] = 1598ns;
slave_timing[1][192+23].t_rxd2[2][1] = 1710ns;

slave_timing[1][192+24].info_corner          = 3;
slave_timing[1][192+24].info_temp__j__       = -40;
slave_timing[1][192+24].info_i__quite_rec__  = 0.040000000;
slave_timing[1][192+24].info_dtr__ib__       = -1;
slave_timing[1][192+24].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+24].info_i__max_slave__  = 0.023000000;
slave_timing[1][192+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][192+24].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+24].t_rxd1[0][1] = 1661ns;
slave_timing[1][192+24].t_rxd1[1][0] = 1648ns;
slave_timing[1][192+24].t_rxd1[0][2] = 1244ns;
slave_timing[1][192+24].t_rxd1[2][0] = 2011ns;
slave_timing[1][192+24].t_rxd2[0][2] = 2000ns;
slave_timing[1][192+24].t_rxd2[2][0] = 1247ns;
slave_timing[1][192+24].t_rxd2[1][2] = 1635ns;
slave_timing[1][192+24].t_rxd2[2][1] = 1655ns;

slave_timing[1][192+25].info_corner          = 3;
slave_timing[1][192+25].info_temp__j__       = -40;
slave_timing[1][192+25].info_i__quite_rec__  = 0.040000000;
slave_timing[1][192+25].info_dtr__ib__       = -1;
slave_timing[1][192+25].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+25].info_i__max_slave__  = 0.025000000;
slave_timing[1][192+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][192+25].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+25].t_rxd1[0][1] = 1594ns;
slave_timing[1][192+25].t_rxd1[1][0] = 1696ns;
slave_timing[1][192+25].t_rxd1[0][2] = 1208ns;
slave_timing[1][192+25].t_rxd1[2][0] = 2046ns;
slave_timing[1][192+25].t_rxd2[0][2] = 1882ns;
slave_timing[1][192+25].t_rxd2[2][0] = 1331ns;
slave_timing[1][192+25].t_rxd2[1][2] = 1463ns;
slave_timing[1][192+25].t_rxd2[2][1] = 1826ns;

slave_timing[1][192+26].info_corner          = 3;
slave_timing[1][192+26].info_temp__j__       = -40;
slave_timing[1][192+26].info_i__quite_rec__  = 0.040000000;
slave_timing[1][192+26].info_dtr__ib__       = 1;
slave_timing[1][192+26].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+26].info_i__max_slave__  = 0.023000000;
slave_timing[1][192+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][192+26].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+26].t_rxd1[0][1] = 1705ns;
slave_timing[1][192+26].t_rxd1[1][0] = 1614ns;
slave_timing[1][192+26].t_rxd1[0][2] = 1266ns;
slave_timing[1][192+26].t_rxd1[2][0] = 1987ns;
slave_timing[1][192+26].t_rxd2[0][2] = 2107ns;
slave_timing[1][192+26].t_rxd2[2][0] = 1181ns;
slave_timing[1][192+26].t_rxd2[1][2] = 1783ns;
slave_timing[1][192+26].t_rxd2[2][1] = 1531ns;

slave_timing[1][192+27].info_corner          = 3;
slave_timing[1][192+27].info_temp__j__       = -40;
slave_timing[1][192+27].info_i__quite_rec__  = 0.040000000;
slave_timing[1][192+27].info_dtr__ib__       = 1;
slave_timing[1][192+27].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+27].info_i__max_slave__  = 0.025000000;
slave_timing[1][192+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][192+27].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+27].t_rxd1[0][1] = 1634ns;
slave_timing[1][192+27].t_rxd1[1][0] = 1662ns;
slave_timing[1][192+27].t_rxd1[0][2] = 1219ns;
slave_timing[1][192+27].t_rxd1[2][0] = 2021ns;
slave_timing[1][192+27].t_rxd2[0][2] = 1947ns;
slave_timing[1][192+27].t_rxd2[2][0] = 1271ns;
slave_timing[1][192+27].t_rxd2[1][2] = 1585ns;
slave_timing[1][192+27].t_rxd2[2][1] = 1704ns;

slave_timing[1][192+28].info_corner          = 3;
slave_timing[1][192+28].info_temp__j__       = -40;
slave_timing[1][192+28].info_i__quite_rec__  = 0.040000000;
slave_timing[1][192+28].info_dtr__ib__       = -1;
slave_timing[1][192+28].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+28].info_i__max_slave__  = 0.023000000;
slave_timing[1][192+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][192+28].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+28].t_rxd1[0][1] = 1701ns;
slave_timing[1][192+28].t_rxd1[1][0] = 1692ns;
slave_timing[1][192+28].t_rxd1[0][2] = 1286ns;
slave_timing[1][192+28].t_rxd1[2][0] = 2051ns;
slave_timing[1][192+28].t_rxd2[0][2] = 2015ns;
slave_timing[1][192+28].t_rxd2[2][0] = 1262ns;
slave_timing[1][192+28].t_rxd2[1][2] = 1651ns;
slave_timing[1][192+28].t_rxd2[2][1] = 1669ns;

slave_timing[1][192+29].info_corner          = 3;
slave_timing[1][192+29].info_temp__j__       = -40;
slave_timing[1][192+29].info_i__quite_rec__  = 0.040000000;
slave_timing[1][192+29].info_dtr__ib__       = -1;
slave_timing[1][192+29].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+29].info_i__max_slave__  = 0.025000000;
slave_timing[1][192+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][192+29].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+29].t_rxd1[0][1] = 1636ns;
slave_timing[1][192+29].t_rxd1[1][0] = 1738ns;
slave_timing[1][192+29].t_rxd1[0][2] = 1247ns;
slave_timing[1][192+29].t_rxd1[2][0] = 2088ns;
slave_timing[1][192+29].t_rxd2[0][2] = 1898ns;
slave_timing[1][192+29].t_rxd2[2][0] = 1347ns;
slave_timing[1][192+29].t_rxd2[1][2] = 1480ns;
slave_timing[1][192+29].t_rxd2[2][1] = 1840ns;

slave_timing[1][192+30].info_corner          = 3;
slave_timing[1][192+30].info_temp__j__       = -40;
slave_timing[1][192+30].info_i__quite_rec__  = 0.040000000;
slave_timing[1][192+30].info_dtr__ib__       = 1;
slave_timing[1][192+30].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+30].info_i__max_slave__  = 0.023000000;
slave_timing[1][192+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][192+30].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+30].t_rxd1[0][1] = 1746ns;
slave_timing[1][192+30].t_rxd1[1][0] = 1656ns;
slave_timing[1][192+30].t_rxd1[0][2] = 1291ns;
slave_timing[1][192+30].t_rxd1[2][0] = 2025ns;
slave_timing[1][192+30].t_rxd2[0][2] = 2120ns;
slave_timing[1][192+30].t_rxd2[2][0] = 1196ns;
slave_timing[1][192+30].t_rxd2[1][2] = 1794ns;
slave_timing[1][192+30].t_rxd2[2][1] = 1543ns;

slave_timing[1][192+31].info_corner          = 3;
slave_timing[1][192+31].info_temp__j__       = -40;
slave_timing[1][192+31].info_i__quite_rec__  = 0.040000000;
slave_timing[1][192+31].info_dtr__ib__       = 1;
slave_timing[1][192+31].info_i__offset_rec__ = 0.000000000;
slave_timing[1][192+31].info_i__max_slave__  = 0.025000000;
slave_timing[1][192+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][192+31].info_r__dsi_bus__    = 5.000;

slave_timing[1][192+31].t_rxd1[0][1] = 1674ns;
slave_timing[1][192+31].t_rxd1[1][0] = 1705ns;
slave_timing[1][192+31].t_rxd1[0][2] = 1266ns;
slave_timing[1][192+31].t_rxd1[2][0] = 2060ns;
slave_timing[1][192+31].t_rxd2[0][2] = 1977ns;
slave_timing[1][192+31].t_rxd2[2][0] = 1286ns;
slave_timing[1][192+31].t_rxd2[1][2] = 1602ns;
slave_timing[1][192+31].t_rxd2[2][1] = 1710ns;

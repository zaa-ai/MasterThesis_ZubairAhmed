my_report_server  = new();
uvm_report_server::set_server( my_report_server );
 

slave_timing[2][224+0].info_corner          = 4;
slave_timing[2][224+0].info_temp__j__       = -40;
slave_timing[2][224+0].info_i__quite_rec__  = 0.006000000;
slave_timing[2][224+0].info_dtr__ib__       = -1;
slave_timing[2][224+0].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+0].info_i__max_slave__  = 0.023000000;
slave_timing[2][224+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][224+0].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+0].t_rxd1[0][1] = 2243ns;
slave_timing[2][224+0].t_rxd1[1][0] = 2200ns;
slave_timing[2][224+0].t_rxd1[0][2] = 1672ns;
slave_timing[2][224+0].t_rxd1[2][0] = 2712ns;
slave_timing[2][224+0].t_rxd2[0][2] = 2684ns;
slave_timing[2][224+0].t_rxd2[2][0] = 1674ns;
slave_timing[2][224+0].t_rxd2[1][2] = 2225ns;
slave_timing[2][224+0].t_rxd2[2][1] = 2198ns;

slave_timing[2][224+1].info_corner          = 4;
slave_timing[2][224+1].info_temp__j__       = -40;
slave_timing[2][224+1].info_i__quite_rec__  = 0.006000000;
slave_timing[2][224+1].info_dtr__ib__       = -1;
slave_timing[2][224+1].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+1].info_i__max_slave__  = 0.025000000;
slave_timing[2][224+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][224+1].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+1].t_rxd1[0][1] = 2137ns;
slave_timing[2][224+1].t_rxd1[1][0] = 2289ns;
slave_timing[2][224+1].t_rxd1[0][2] = 1640ns;
slave_timing[2][224+1].t_rxd1[2][0] = 2759ns;
slave_timing[2][224+1].t_rxd2[0][2] = 2552ns;
slave_timing[2][224+1].t_rxd2[2][0] = 1789ns;
slave_timing[2][224+1].t_rxd2[1][2] = 2002ns;
slave_timing[2][224+1].t_rxd2[2][1] = 2393ns;

slave_timing[2][224+2].info_corner          = 4;
slave_timing[2][224+2].info_temp__j__       = -40;
slave_timing[2][224+2].info_i__quite_rec__  = 0.006000000;
slave_timing[2][224+2].info_dtr__ib__       = 1;
slave_timing[2][224+2].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+2].info_i__max_slave__  = 0.023000000;
slave_timing[2][224+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][224+2].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+2].t_rxd1[0][1] = 2290ns;
slave_timing[2][224+2].t_rxd1[1][0] = 2183ns;
slave_timing[2][224+2].t_rxd1[0][2] = 1714ns;
slave_timing[2][224+2].t_rxd1[2][0] = 2687ns;
slave_timing[2][224+2].t_rxd2[0][2] = 2832ns;
slave_timing[2][224+2].t_rxd2[2][0] = 1586ns;
slave_timing[2][224+2].t_rxd2[1][2] = 2397ns;
slave_timing[2][224+2].t_rxd2[2][1] = 2049ns;

slave_timing[2][224+3].info_corner          = 4;
slave_timing[2][224+3].info_temp__j__       = -40;
slave_timing[2][224+3].info_i__quite_rec__  = 0.006000000;
slave_timing[2][224+3].info_dtr__ib__       = 1;
slave_timing[2][224+3].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+3].info_i__max_slave__  = 0.025000000;
slave_timing[2][224+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][224+3].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+3].t_rxd1[0][1] = 2197ns;
slave_timing[2][224+3].t_rxd1[1][0] = 2251ns;
slave_timing[2][224+3].t_rxd1[0][2] = 1663ns;
slave_timing[2][224+3].t_rxd1[2][0] = 2732ns;
slave_timing[2][224+3].t_rxd2[0][2] = 2642ns;
slave_timing[2][224+3].t_rxd2[2][0] = 1719ns;
slave_timing[2][224+3].t_rxd2[1][2] = 2139ns;
slave_timing[2][224+3].t_rxd2[2][1] = 2249ns;

slave_timing[2][224+4].info_corner          = 4;
slave_timing[2][224+4].info_temp__j__       = -40;
slave_timing[2][224+4].info_i__quite_rec__  = 0.006000000;
slave_timing[2][224+4].info_dtr__ib__       = -1;
slave_timing[2][224+4].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+4].info_i__max_slave__  = 0.023000000;
slave_timing[2][224+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][224+4].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+4].t_rxd1[0][1] = 2323ns;
slave_timing[2][224+4].t_rxd1[1][0] = 2284ns;
slave_timing[2][224+4].t_rxd1[0][2] = 1733ns;
slave_timing[2][224+4].t_rxd1[2][0] = 2778ns;
slave_timing[2][224+4].t_rxd2[0][2] = 2700ns;
slave_timing[2][224+4].t_rxd2[2][0] = 1687ns;
slave_timing[2][224+4].t_rxd2[1][2] = 2249ns;
slave_timing[2][224+4].t_rxd2[2][1] = 2215ns;

slave_timing[2][224+5].info_corner          = 4;
slave_timing[2][224+5].info_temp__j__       = -40;
slave_timing[2][224+5].info_i__quite_rec__  = 0.006000000;
slave_timing[2][224+5].info_dtr__ib__       = -1;
slave_timing[2][224+5].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+5].info_i__max_slave__  = 0.025000000;
slave_timing[2][224+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][224+5].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+5].t_rxd1[0][1] = 2231ns;
slave_timing[2][224+5].t_rxd1[1][0] = 2357ns;
slave_timing[2][224+5].t_rxd1[0][2] = 1703ns;
slave_timing[2][224+5].t_rxd1[2][0] = 2822ns;
slave_timing[2][224+5].t_rxd2[0][2] = 2568ns;
slave_timing[2][224+5].t_rxd2[2][0] = 1801ns;
slave_timing[2][224+5].t_rxd2[1][2] = 2011ns;
slave_timing[2][224+5].t_rxd2[2][1] = 2439ns;

slave_timing[2][224+6].info_corner          = 4;
slave_timing[2][224+6].info_temp__j__       = -40;
slave_timing[2][224+6].info_i__quite_rec__  = 0.006000000;
slave_timing[2][224+6].info_dtr__ib__       = 1;
slave_timing[2][224+6].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+6].info_i__max_slave__  = 0.023000000;
slave_timing[2][224+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][224+6].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+6].t_rxd1[0][1] = 2368ns;
slave_timing[2][224+6].t_rxd1[1][0] = 2251ns;
slave_timing[2][224+6].t_rxd1[0][2] = 1776ns;
slave_timing[2][224+6].t_rxd1[2][0] = 2748ns;
slave_timing[2][224+6].t_rxd2[0][2] = 2837ns;
slave_timing[2][224+6].t_rxd2[2][0] = 1598ns;
slave_timing[2][224+6].t_rxd2[1][2] = 2416ns;
slave_timing[2][224+6].t_rxd2[2][1] = 2060ns;

slave_timing[2][224+7].info_corner          = 4;
slave_timing[2][224+7].info_temp__j__       = -40;
slave_timing[2][224+7].info_i__quite_rec__  = 0.006000000;
slave_timing[2][224+7].info_dtr__ib__       = 1;
slave_timing[2][224+7].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+7].info_i__max_slave__  = 0.025000000;
slave_timing[2][224+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][224+7].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+7].t_rxd1[0][1] = 2268ns;
slave_timing[2][224+7].t_rxd1[1][0] = 2317ns;
slave_timing[2][224+7].t_rxd1[0][2] = 1722ns;
slave_timing[2][224+7].t_rxd1[2][0] = 2787ns;
slave_timing[2][224+7].t_rxd2[0][2] = 2664ns;
slave_timing[2][224+7].t_rxd2[2][0] = 1729ns;
slave_timing[2][224+7].t_rxd2[1][2] = 2148ns;
slave_timing[2][224+7].t_rxd2[2][1] = 2298ns;

slave_timing[2][224+8].info_corner          = 4;
slave_timing[2][224+8].info_temp__j__       = -40;
slave_timing[2][224+8].info_i__quite_rec__  = 0.003000000;
slave_timing[2][224+8].info_dtr__ib__       = -1;
slave_timing[2][224+8].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+8].info_i__max_slave__  = 0.023000000;
slave_timing[2][224+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][224+8].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+8].t_rxd1[0][1] = 2225ns;
slave_timing[2][224+8].t_rxd1[1][0] = 2240ns;
slave_timing[2][224+8].t_rxd1[0][2] = 1674ns;
slave_timing[2][224+8].t_rxd1[2][0] = 2726ns;
slave_timing[2][224+8].t_rxd2[0][2] = 2695ns;
slave_timing[2][224+8].t_rxd2[2][0] = 1679ns;
slave_timing[2][224+8].t_rxd2[1][2] = 2200ns;
slave_timing[2][224+8].t_rxd2[2][1] = 2181ns;

slave_timing[2][224+9].info_corner          = 4;
slave_timing[2][224+9].info_temp__j__       = -40;
slave_timing[2][224+9].info_i__quite_rec__  = 0.003000000;
slave_timing[2][224+9].info_dtr__ib__       = -1;
slave_timing[2][224+9].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+9].info_i__max_slave__  = 0.025000000;
slave_timing[2][224+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][224+9].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+9].t_rxd1[0][1] = 2139ns;
slave_timing[2][224+9].t_rxd1[1][0] = 2296ns;
slave_timing[2][224+9].t_rxd1[0][2] = 1629ns;
slave_timing[2][224+9].t_rxd1[2][0] = 2768ns;
slave_timing[2][224+9].t_rxd2[0][2] = 2544ns;
slave_timing[2][224+9].t_rxd2[2][0] = 1795ns;
slave_timing[2][224+9].t_rxd2[1][2] = 1976ns;
slave_timing[2][224+9].t_rxd2[2][1] = 2442ns;

slave_timing[2][224+10].info_corner          = 4;
slave_timing[2][224+10].info_temp__j__       = -40;
slave_timing[2][224+10].info_i__quite_rec__  = 0.003000000;
slave_timing[2][224+10].info_dtr__ib__       = 1;
slave_timing[2][224+10].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+10].info_i__max_slave__  = 0.023000000;
slave_timing[2][224+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][224+10].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+10].t_rxd1[0][1] = 2277ns;
slave_timing[2][224+10].t_rxd1[1][0] = 2191ns;
slave_timing[2][224+10].t_rxd1[0][2] = 1710ns;
slave_timing[2][224+10].t_rxd1[2][0] = 2690ns;
slave_timing[2][224+10].t_rxd2[0][2] = 2815ns;
slave_timing[2][224+10].t_rxd2[2][0] = 1591ns;
slave_timing[2][224+10].t_rxd2[1][2] = 2390ns;
slave_timing[2][224+10].t_rxd2[2][1] = 2055ns;

slave_timing[2][224+11].info_corner          = 4;
slave_timing[2][224+11].info_temp__j__       = -40;
slave_timing[2][224+11].info_i__quite_rec__  = 0.003000000;
slave_timing[2][224+11].info_dtr__ib__       = 1;
slave_timing[2][224+11].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+11].info_i__max_slave__  = 0.025000000;
slave_timing[2][224+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][224+11].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+11].t_rxd1[0][1] = 2190ns;
slave_timing[2][224+11].t_rxd1[1][0] = 2252ns;
slave_timing[2][224+11].t_rxd1[0][2] = 1657ns;
slave_timing[2][224+11].t_rxd1[2][0] = 2738ns;
slave_timing[2][224+11].t_rxd2[0][2] = 2638ns;
slave_timing[2][224+11].t_rxd2[2][0] = 1720ns;
slave_timing[2][224+11].t_rxd2[1][2] = 2127ns;
slave_timing[2][224+11].t_rxd2[2][1] = 2291ns;

slave_timing[2][224+12].info_corner          = 4;
slave_timing[2][224+12].info_temp__j__       = -40;
slave_timing[2][224+12].info_i__quite_rec__  = 0.003000000;
slave_timing[2][224+12].info_dtr__ib__       = -1;
slave_timing[2][224+12].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+12].info_i__max_slave__  = 0.023000000;
slave_timing[2][224+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][224+12].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+12].t_rxd1[0][1] = 2299ns;
slave_timing[2][224+12].t_rxd1[1][0] = 2309ns;
slave_timing[2][224+12].t_rxd1[0][2] = 1747ns;
slave_timing[2][224+12].t_rxd1[2][0] = 2791ns;
slave_timing[2][224+12].t_rxd2[0][2] = 2712ns;
slave_timing[2][224+12].t_rxd2[2][0] = 1692ns;
slave_timing[2][224+12].t_rxd2[1][2] = 2227ns;
slave_timing[2][224+12].t_rxd2[2][1] = 2221ns;

slave_timing[2][224+13].info_corner          = 4;
slave_timing[2][224+13].info_temp__j__       = -40;
slave_timing[2][224+13].info_i__quite_rec__  = 0.003000000;
slave_timing[2][224+13].info_dtr__ib__       = -1;
slave_timing[2][224+13].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+13].info_i__max_slave__  = 0.025000000;
slave_timing[2][224+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][224+13].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+13].t_rxd1[0][1] = 2221ns;
slave_timing[2][224+13].t_rxd1[1][0] = 2378ns;
slave_timing[2][224+13].t_rxd1[0][2] = 1697ns;
slave_timing[2][224+13].t_rxd1[2][0] = 2838ns;
slave_timing[2][224+13].t_rxd2[0][2] = 2558ns;
slave_timing[2][224+13].t_rxd2[2][0] = 1808ns;
slave_timing[2][224+13].t_rxd2[1][2] = 1994ns;
slave_timing[2][224+13].t_rxd2[2][1] = 2450ns;

slave_timing[2][224+14].info_corner          = 4;
slave_timing[2][224+14].info_temp__j__       = -40;
slave_timing[2][224+14].info_i__quite_rec__  = 0.003000000;
slave_timing[2][224+14].info_dtr__ib__       = 1;
slave_timing[2][224+14].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+14].info_i__max_slave__  = 0.023000000;
slave_timing[2][224+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][224+14].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+14].t_rxd1[0][1] = 2351ns;
slave_timing[2][224+14].t_rxd1[1][0] = 2265ns;
slave_timing[2][224+14].t_rxd1[0][2] = 1770ns;
slave_timing[2][224+14].t_rxd1[2][0] = 2756ns;
slave_timing[2][224+14].t_rxd2[0][2] = 2829ns;
slave_timing[2][224+14].t_rxd2[2][0] = 1603ns;
slave_timing[2][224+14].t_rxd2[1][2] = 2400ns;
slave_timing[2][224+14].t_rxd2[2][1] = 2060ns;

slave_timing[2][224+15].info_corner          = 4;
slave_timing[2][224+15].info_temp__j__       = -40;
slave_timing[2][224+15].info_i__quite_rec__  = 0.003000000;
slave_timing[2][224+15].info_dtr__ib__       = 1;
slave_timing[2][224+15].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+15].info_i__max_slave__  = 0.025000000;
slave_timing[2][224+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][224+15].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+15].t_rxd1[0][1] = 2264ns;
slave_timing[2][224+15].t_rxd1[1][0] = 2322ns;
slave_timing[2][224+15].t_rxd1[0][2] = 1719ns;
slave_timing[2][224+15].t_rxd1[2][0] = 2799ns;
slave_timing[2][224+15].t_rxd2[0][2] = 2650ns;
slave_timing[2][224+15].t_rxd2[2][0] = 1735ns;
slave_timing[2][224+15].t_rxd2[1][2] = 2138ns;
slave_timing[2][224+15].t_rxd2[2][1] = 2304ns;

slave_timing[2][224+16].info_corner          = 4;
slave_timing[2][224+16].info_temp__j__       = -40;
slave_timing[2][224+16].info_i__quite_rec__  = 0.000000000;
slave_timing[2][224+16].info_dtr__ib__       = -1;
slave_timing[2][224+16].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+16].info_i__max_slave__  = 0.023000000;
slave_timing[2][224+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][224+16].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+16].t_rxd1[0][1] = 2247ns;
slave_timing[2][224+16].t_rxd1[1][0] = 2224ns;
slave_timing[2][224+16].t_rxd1[0][2] = 1673ns;
slave_timing[2][224+16].t_rxd1[2][0] = 2714ns;
slave_timing[2][224+16].t_rxd2[0][2] = 2686ns;
slave_timing[2][224+16].t_rxd2[2][0] = 1675ns;
slave_timing[2][224+16].t_rxd2[1][2] = 2229ns;
slave_timing[2][224+16].t_rxd2[2][1] = 2209ns;

slave_timing[2][224+17].info_corner          = 4;
slave_timing[2][224+17].info_temp__j__       = -40;
slave_timing[2][224+17].info_i__quite_rec__  = 0.000000000;
slave_timing[2][224+17].info_dtr__ib__       = -1;
slave_timing[2][224+17].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+17].info_i__max_slave__  = 0.025000000;
slave_timing[2][224+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][224+17].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+17].t_rxd1[0][1] = 2160ns;
slave_timing[2][224+17].t_rxd1[1][0] = 2290ns;
slave_timing[2][224+17].t_rxd1[0][2] = 1623ns;
slave_timing[2][224+17].t_rxd1[2][0] = 2784ns;
slave_timing[2][224+17].t_rxd2[0][2] = 2535ns;
slave_timing[2][224+17].t_rxd2[2][0] = 1807ns;
slave_timing[2][224+17].t_rxd2[1][2] = 1994ns;
slave_timing[2][224+17].t_rxd2[2][1] = 2437ns;

slave_timing[2][224+18].info_corner          = 4;
slave_timing[2][224+18].info_temp__j__       = -40;
slave_timing[2][224+18].info_i__quite_rec__  = 0.000000000;
slave_timing[2][224+18].info_dtr__ib__       = 1;
slave_timing[2][224+18].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+18].info_i__max_slave__  = 0.023000000;
slave_timing[2][224+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][224+18].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+18].t_rxd1[0][1] = 2276ns;
slave_timing[2][224+18].t_rxd1[1][0] = 2208ns;
slave_timing[2][224+18].t_rxd1[0][2] = 1705ns;
slave_timing[2][224+18].t_rxd1[2][0] = 2701ns;
slave_timing[2][224+18].t_rxd2[0][2] = 2804ns;
slave_timing[2][224+18].t_rxd2[2][0] = 1592ns;
slave_timing[2][224+18].t_rxd2[1][2] = 2408ns;
slave_timing[2][224+18].t_rxd2[2][1] = 2038ns;

slave_timing[2][224+19].info_corner          = 4;
slave_timing[2][224+19].info_temp__j__       = -40;
slave_timing[2][224+19].info_i__quite_rec__  = 0.000000000;
slave_timing[2][224+19].info_dtr__ib__       = 1;
slave_timing[2][224+19].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+19].info_i__max_slave__  = 0.025000000;
slave_timing[2][224+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][224+19].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+19].t_rxd1[0][1] = 2181ns;
slave_timing[2][224+19].t_rxd1[1][0] = 2278ns;
slave_timing[2][224+19].t_rxd1[0][2] = 1655ns;
slave_timing[2][224+19].t_rxd1[2][0] = 2755ns;
slave_timing[2][224+19].t_rxd2[0][2] = 2632ns;
slave_timing[2][224+19].t_rxd2[2][0] = 1728ns;
slave_timing[2][224+19].t_rxd2[1][2] = 2118ns;
slave_timing[2][224+19].t_rxd2[2][1] = 2300ns;

slave_timing[2][224+20].info_corner          = 4;
slave_timing[2][224+20].info_temp__j__       = -40;
slave_timing[2][224+20].info_i__quite_rec__  = 0.000000000;
slave_timing[2][224+20].info_dtr__ib__       = -1;
slave_timing[2][224+20].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+20].info_i__max_slave__  = 0.023000000;
slave_timing[2][224+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][224+20].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+20].t_rxd1[0][1] = 2323ns;
slave_timing[2][224+20].t_rxd1[1][0] = 2286ns;
slave_timing[2][224+20].t_rxd1[0][2] = 1739ns;
slave_timing[2][224+20].t_rxd1[2][0] = 2782ns;
slave_timing[2][224+20].t_rxd2[0][2] = 2698ns;
slave_timing[2][224+20].t_rxd2[2][0] = 1686ns;
slave_timing[2][224+20].t_rxd2[1][2] = 2240ns;
slave_timing[2][224+20].t_rxd2[2][1] = 2205ns;

slave_timing[2][224+21].info_corner          = 4;
slave_timing[2][224+21].info_temp__j__       = -40;
slave_timing[2][224+21].info_i__quite_rec__  = 0.000000000;
slave_timing[2][224+21].info_dtr__ib__       = -1;
slave_timing[2][224+21].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+21].info_i__max_slave__  = 0.025000000;
slave_timing[2][224+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][224+21].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+21].t_rxd1[0][1] = 2208ns;
slave_timing[2][224+21].t_rxd1[1][0] = 2389ns;
slave_timing[2][224+21].t_rxd1[0][2] = 1691ns;
slave_timing[2][224+21].t_rxd1[2][0] = 2845ns;
slave_timing[2][224+21].t_rxd2[0][2] = 2550ns;
slave_timing[2][224+21].t_rxd2[2][0] = 1819ns;
slave_timing[2][224+21].t_rxd2[1][2] = 2011ns;
slave_timing[2][224+21].t_rxd2[2][1] = 2442ns;

slave_timing[2][224+22].info_corner          = 4;
slave_timing[2][224+22].info_temp__j__       = -40;
slave_timing[2][224+22].info_i__quite_rec__  = 0.000000000;
slave_timing[2][224+22].info_dtr__ib__       = 1;
slave_timing[2][224+22].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+22].info_i__max_slave__  = 0.023000000;
slave_timing[2][224+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][224+22].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+22].t_rxd1[0][1] = 2347ns;
slave_timing[2][224+22].t_rxd1[1][0] = 2268ns;
slave_timing[2][224+22].t_rxd1[0][2] = 1765ns;
slave_timing[2][224+22].t_rxd1[2][0] = 2766ns;
slave_timing[2][224+22].t_rxd2[0][2] = 2816ns;
slave_timing[2][224+22].t_rxd2[2][0] = 1609ns;
slave_timing[2][224+22].t_rxd2[1][2] = 2424ns;
slave_timing[2][224+22].t_rxd2[2][1] = 2050ns;

slave_timing[2][224+23].info_corner          = 4;
slave_timing[2][224+23].info_temp__j__       = -40;
slave_timing[2][224+23].info_i__quite_rec__  = 0.000000000;
slave_timing[2][224+23].info_dtr__ib__       = 1;
slave_timing[2][224+23].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+23].info_i__max_slave__  = 0.025000000;
slave_timing[2][224+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][224+23].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+23].t_rxd1[0][1] = 2251ns;
slave_timing[2][224+23].t_rxd1[1][0] = 2340ns;
slave_timing[2][224+23].t_rxd1[0][2] = 1713ns;
slave_timing[2][224+23].t_rxd1[2][0] = 2810ns;
slave_timing[2][224+23].t_rxd2[0][2] = 2641ns;
slave_timing[2][224+23].t_rxd2[2][0] = 1739ns;
slave_timing[2][224+23].t_rxd2[1][2] = 2134ns;
slave_timing[2][224+23].t_rxd2[2][1] = 2315ns;

slave_timing[2][224+24].info_corner          = 4;
slave_timing[2][224+24].info_temp__j__       = -40;
slave_timing[2][224+24].info_i__quite_rec__  = 0.040000000;
slave_timing[2][224+24].info_dtr__ib__       = -1;
slave_timing[2][224+24].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+24].info_i__max_slave__  = 0.023000000;
slave_timing[2][224+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][224+24].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+24].t_rxd1[0][1] = 2199ns;
slave_timing[2][224+24].t_rxd1[1][0] = 2238ns;
slave_timing[2][224+24].t_rxd1[0][2] = 1666ns;
slave_timing[2][224+24].t_rxd1[2][0] = 2726ns;
slave_timing[2][224+24].t_rxd2[0][2] = 2689ns;
slave_timing[2][224+24].t_rxd2[2][0] = 1678ns;
slave_timing[2][224+24].t_rxd2[1][2] = 2200ns;
slave_timing[2][224+24].t_rxd2[2][1] = 2225ns;

slave_timing[2][224+25].info_corner          = 4;
slave_timing[2][224+25].info_temp__j__       = -40;
slave_timing[2][224+25].info_i__quite_rec__  = 0.040000000;
slave_timing[2][224+25].info_dtr__ib__       = -1;
slave_timing[2][224+25].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+25].info_i__max_slave__  = 0.025000000;
slave_timing[2][224+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][224+25].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+25].t_rxd1[0][1] = 2122ns;
slave_timing[2][224+25].t_rxd1[1][0] = 2300ns;
slave_timing[2][224+25].t_rxd1[0][2] = 1615ns;
slave_timing[2][224+25].t_rxd1[2][0] = 2763ns;
slave_timing[2][224+25].t_rxd2[0][2] = 2534ns;
slave_timing[2][224+25].t_rxd2[2][0] = 1798ns;
slave_timing[2][224+25].t_rxd2[1][2] = 1976ns;
slave_timing[2][224+25].t_rxd2[2][1] = 2426ns;

slave_timing[2][224+26].info_corner          = 4;
slave_timing[2][224+26].info_temp__j__       = -40;
slave_timing[2][224+26].info_i__quite_rec__  = 0.040000000;
slave_timing[2][224+26].info_dtr__ib__       = 1;
slave_timing[2][224+26].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+26].info_i__max_slave__  = 0.023000000;
slave_timing[2][224+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][224+26].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+26].t_rxd1[0][1] = 2276ns;
slave_timing[2][224+26].t_rxd1[1][0] = 2167ns;
slave_timing[2][224+26].t_rxd1[0][2] = 1704ns;
slave_timing[2][224+26].t_rxd1[2][0] = 2679ns;
slave_timing[2][224+26].t_rxd2[0][2] = 2819ns;
slave_timing[2][224+26].t_rxd2[2][0] = 1584ns;
slave_timing[2][224+26].t_rxd2[1][2] = 2406ns;
slave_timing[2][224+26].t_rxd2[2][1] = 2055ns;

slave_timing[2][224+27].info_corner          = 4;
slave_timing[2][224+27].info_temp__j__       = -40;
slave_timing[2][224+27].info_i__quite_rec__  = 0.040000000;
slave_timing[2][224+27].info_dtr__ib__       = 1;
slave_timing[2][224+27].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+27].info_i__max_slave__  = 0.025000000;
slave_timing[2][224+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][224+27].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+27].t_rxd1[0][1] = 2185ns;
slave_timing[2][224+27].t_rxd1[1][0] = 2246ns;
slave_timing[2][224+27].t_rxd1[0][2] = 1651ns;
slave_timing[2][224+27].t_rxd1[2][0] = 2726ns;
slave_timing[2][224+27].t_rxd2[0][2] = 2639ns;
slave_timing[2][224+27].t_rxd2[2][0] = 1710ns;
slave_timing[2][224+27].t_rxd2[1][2] = 2129ns;
slave_timing[2][224+27].t_rxd2[2][1] = 2288ns;

slave_timing[2][224+28].info_corner          = 4;
slave_timing[2][224+28].info_temp__j__       = -40;
slave_timing[2][224+28].info_i__quite_rec__  = 0.040000000;
slave_timing[2][224+28].info_dtr__ib__       = -1;
slave_timing[2][224+28].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+28].info_i__max_slave__  = 0.023000000;
slave_timing[2][224+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][224+28].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+28].t_rxd1[0][1] = 2240ns;
slave_timing[2][224+28].t_rxd1[1][0] = 2269ns;
slave_timing[2][224+28].t_rxd1[0][2] = 1701ns;
slave_timing[2][224+28].t_rxd1[2][0] = 2754ns;
slave_timing[2][224+28].t_rxd2[0][2] = 2700ns;
slave_timing[2][224+28].t_rxd2[2][0] = 1698ns;
slave_timing[2][224+28].t_rxd2[1][2] = 2224ns;
slave_timing[2][224+28].t_rxd2[2][1] = 2232ns;

slave_timing[2][224+29].info_corner          = 4;
slave_timing[2][224+29].info_temp__j__       = -40;
slave_timing[2][224+29].info_i__quite_rec__  = 0.040000000;
slave_timing[2][224+29].info_dtr__ib__       = -1;
slave_timing[2][224+29].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+29].info_i__max_slave__  = 0.025000000;
slave_timing[2][224+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][224+29].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+29].t_rxd1[0][1] = 2162ns;
slave_timing[2][224+29].t_rxd1[1][0] = 2335ns;
slave_timing[2][224+29].t_rxd1[0][2] = 1650ns;
slave_timing[2][224+29].t_rxd1[2][0] = 2798ns;
slave_timing[2][224+29].t_rxd2[0][2] = 2557ns;
slave_timing[2][224+29].t_rxd2[2][0] = 1814ns;
slave_timing[2][224+29].t_rxd2[1][2] = 1988ns;
slave_timing[2][224+29].t_rxd2[2][1] = 2465ns;

slave_timing[2][224+30].info_corner          = 4;
slave_timing[2][224+30].info_temp__j__       = -40;
slave_timing[2][224+30].info_i__quite_rec__  = 0.040000000;
slave_timing[2][224+30].info_dtr__ib__       = 1;
slave_timing[2][224+30].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+30].info_i__max_slave__  = 0.023000000;
slave_timing[2][224+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][224+30].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+30].t_rxd1[0][1] = 2311ns;
slave_timing[2][224+30].t_rxd1[1][0] = 2212ns;
slave_timing[2][224+30].t_rxd1[0][2] = 1733ns;
slave_timing[2][224+30].t_rxd1[2][0] = 2711ns;
slave_timing[2][224+30].t_rxd2[0][2] = 2826ns;
slave_timing[2][224+30].t_rxd2[2][0] = 1600ns;
slave_timing[2][224+30].t_rxd2[1][2] = 2407ns;
slave_timing[2][224+30].t_rxd2[2][1] = 2072ns;

slave_timing[2][224+31].info_corner          = 4;
slave_timing[2][224+31].info_temp__j__       = -40;
slave_timing[2][224+31].info_i__quite_rec__  = 0.040000000;
slave_timing[2][224+31].info_dtr__ib__       = 1;
slave_timing[2][224+31].info_i__offset_rec__ = 0.000000000;
slave_timing[2][224+31].info_i__max_slave__  = 0.025000000;
slave_timing[2][224+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][224+31].info_r__dsi_bus__    = 5.000;

slave_timing[2][224+31].t_rxd1[0][1] = 2212ns;
slave_timing[2][224+31].t_rxd1[1][0] = 2285ns;
slave_timing[2][224+31].t_rxd1[0][2] = 1682ns;
slave_timing[2][224+31].t_rxd1[2][0] = 2756ns;
slave_timing[2][224+31].t_rxd2[0][2] = 2655ns;
slave_timing[2][224+31].t_rxd2[2][0] = 1725ns;
slave_timing[2][224+31].t_rxd2[1][2] = 2156ns;
slave_timing[2][224+31].t_rxd2[2][1] = 2302ns;

`include "dsi3_master_subscriber.svh"

/* ###   interface instances   ###################################################### */

time_base_registers_TRIM_OSC_if time_base_registers_TRIM_OSC (); 
time_base_registers_TRIM_OSC_TCF_if time_base_registers_TRIM_OSC_TCF (); 
time_base_registers_CLKREF_CONF_if time_base_registers_CLKREF_CONF (); 
time_base_registers_TB_CNT_if time_base_registers_TB_CNT (); 



slave_timing[0][128+0].info_corner          = 1;
slave_timing[0][128+0].info_temp__j__       = -40;
slave_timing[0][128+0].info_i__quite_rec__  = 0.006000000;
slave_timing[0][128+0].info_dtr__ib__       = -1;
slave_timing[0][128+0].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+0].info_i__max_slave__  = 0.023000000;
slave_timing[0][128+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][128+0].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+0].t_rxd1[0][1] = 1059ns;
slave_timing[0][128+0].t_rxd1[1][0] = 1089ns;
slave_timing[0][128+0].t_rxd1[0][2] = 778ns;
slave_timing[0][128+0].t_rxd1[2][0] = 1360ns;
slave_timing[0][128+0].t_rxd2[0][2] = 1296ns;
slave_timing[0][128+0].t_rxd2[2][0] = 800ns;
slave_timing[0][128+0].t_rxd2[1][2] = 1036ns;
slave_timing[0][128+0].t_rxd2[2][1] = 1074ns;

slave_timing[0][128+1].info_corner          = 1;
slave_timing[0][128+1].info_temp__j__       = -40;
slave_timing[0][128+1].info_i__quite_rec__  = 0.006000000;
slave_timing[0][128+1].info_dtr__ib__       = -1;
slave_timing[0][128+1].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+1].info_i__max_slave__  = 0.025000000;
slave_timing[0][128+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][128+1].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+1].t_rxd1[0][1] = 1015ns;
slave_timing[0][128+1].t_rxd1[1][0] = 1124ns;
slave_timing[0][128+1].t_rxd1[0][2] = 765ns;
slave_timing[0][128+1].t_rxd1[2][0] = 1386ns;
slave_timing[0][128+1].t_rxd2[0][2] = 1218ns;
slave_timing[0][128+1].t_rxd2[2][0] = 850ns;
slave_timing[0][128+1].t_rxd2[1][2] = 917ns;
slave_timing[0][128+1].t_rxd2[2][1] = 1202ns;

slave_timing[0][128+2].info_corner          = 1;
slave_timing[0][128+2].info_temp__j__       = -40;
slave_timing[0][128+2].info_i__quite_rec__  = 0.006000000;
slave_timing[0][128+2].info_dtr__ib__       = 1;
slave_timing[0][128+2].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+2].info_i__max_slave__  = 0.023000000;
slave_timing[0][128+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][128+2].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+2].t_rxd1[0][1] = 1106ns;
slave_timing[0][128+2].t_rxd1[1][0] = 1053ns;
slave_timing[0][128+2].t_rxd1[0][2] = 806ns;
slave_timing[0][128+2].t_rxd1[2][0] = 1329ns;
slave_timing[0][128+2].t_rxd2[0][2] = 1416ns;
slave_timing[0][128+2].t_rxd2[2][0] = 744ns;
slave_timing[0][128+2].t_rxd2[1][2] = 1162ns;
slave_timing[0][128+2].t_rxd2[2][1] = 973ns;

slave_timing[0][128+3].info_corner          = 1;
slave_timing[0][128+3].info_temp__j__       = -40;
slave_timing[0][128+3].info_i__quite_rec__  = 0.006000000;
slave_timing[0][128+3].info_dtr__ib__       = 1;
slave_timing[0][128+3].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+3].info_i__max_slave__  = 0.025000000;
slave_timing[0][128+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][128+3].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+3].t_rxd1[0][1] = 1057ns;
slave_timing[0][128+3].t_rxd1[1][0] = 1090ns;
slave_timing[0][128+3].t_rxd1[0][2] = 785ns;
slave_timing[0][128+3].t_rxd1[2][0] = 1359ns;
slave_timing[0][128+3].t_rxd2[0][2] = 1296ns;
slave_timing[0][128+3].t_rxd2[2][0] = 805ns;
slave_timing[0][128+3].t_rxd2[1][2] = 1018ns;
slave_timing[0][128+3].t_rxd2[2][1] = 1091ns;

slave_timing[0][128+4].info_corner          = 1;
slave_timing[0][128+4].info_temp__j__       = -40;
slave_timing[0][128+4].info_i__quite_rec__  = 0.006000000;
slave_timing[0][128+4].info_dtr__ib__       = -1;
slave_timing[0][128+4].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+4].info_i__max_slave__  = 0.023000000;
slave_timing[0][128+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][128+4].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+4].t_rxd1[0][1] = 1137ns;
slave_timing[0][128+4].t_rxd1[1][0] = 1161ns;
slave_timing[0][128+4].t_rxd1[0][2] = 848ns;
slave_timing[0][128+4].t_rxd1[2][0] = 1425ns;
slave_timing[0][128+4].t_rxd2[0][2] = 1333ns;
slave_timing[0][128+4].t_rxd2[2][0] = 819ns;
slave_timing[0][128+4].t_rxd2[1][2] = 1051ns;
slave_timing[0][128+4].t_rxd2[2][1] = 1088ns;

slave_timing[0][128+5].info_corner          = 1;
slave_timing[0][128+5].info_temp__j__       = -40;
slave_timing[0][128+5].info_i__quite_rec__  = 0.006000000;
slave_timing[0][128+5].info_dtr__ib__       = -1;
slave_timing[0][128+5].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+5].info_i__max_slave__  = 0.025000000;
slave_timing[0][128+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][128+5].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+5].t_rxd1[0][1] = 1091ns;
slave_timing[0][128+5].t_rxd1[1][0] = 1195ns;
slave_timing[0][128+5].t_rxd1[0][2] = 825ns;
slave_timing[0][128+5].t_rxd1[2][0] = 1453ns;
slave_timing[0][128+5].t_rxd2[0][2] = 1242ns;
slave_timing[0][128+5].t_rxd2[2][0] = 872ns;
slave_timing[0][128+5].t_rxd2[1][2] = 934ns;
slave_timing[0][128+5].t_rxd2[2][1] = 1217ns;

slave_timing[0][128+6].info_corner          = 1;
slave_timing[0][128+6].info_temp__j__       = -40;
slave_timing[0][128+6].info_i__quite_rec__  = 0.006000000;
slave_timing[0][128+6].info_dtr__ib__       = 1;
slave_timing[0][128+6].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+6].info_i__max_slave__  = 0.023000000;
slave_timing[0][128+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][128+6].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+6].t_rxd1[0][1] = 1186ns;
slave_timing[0][128+6].t_rxd1[1][0] = 1125ns;
slave_timing[0][128+6].t_rxd1[0][2] = 871ns;
slave_timing[0][128+6].t_rxd1[2][0] = 1398ns;
slave_timing[0][128+6].t_rxd2[0][2] = 1439ns;
slave_timing[0][128+6].t_rxd2[2][0] = 767ns;
slave_timing[0][128+6].t_rxd2[1][2] = 1174ns;
slave_timing[0][128+6].t_rxd2[2][1] = 987ns;

slave_timing[0][128+7].info_corner          = 1;
slave_timing[0][128+7].info_temp__j__       = -40;
slave_timing[0][128+7].info_i__quite_rec__  = 0.006000000;
slave_timing[0][128+7].info_dtr__ib__       = 1;
slave_timing[0][128+7].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+7].info_i__max_slave__  = 0.025000000;
slave_timing[0][128+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][128+7].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+7].t_rxd1[0][1] = 1133ns;
slave_timing[0][128+7].t_rxd1[1][0] = 1162ns;
slave_timing[0][128+7].t_rxd1[0][2] = 845ns;
slave_timing[0][128+7].t_rxd1[2][0] = 1424ns;
slave_timing[0][128+7].t_rxd2[0][2] = 1318ns;
slave_timing[0][128+7].t_rxd2[2][0] = 822ns;
slave_timing[0][128+7].t_rxd2[1][2] = 1035ns;
slave_timing[0][128+7].t_rxd2[2][1] = 1086ns;

slave_timing[0][128+8].info_corner          = 1;
slave_timing[0][128+8].info_temp__j__       = -40;
slave_timing[0][128+8].info_i__quite_rec__  = 0.003000000;
slave_timing[0][128+8].info_dtr__ib__       = -1;
slave_timing[0][128+8].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+8].info_i__max_slave__  = 0.023000000;
slave_timing[0][128+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][128+8].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+8].t_rxd1[0][1] = 1072ns;
slave_timing[0][128+8].t_rxd1[1][0] = 1076ns;
slave_timing[0][128+8].t_rxd1[0][2] = 792ns;
slave_timing[0][128+8].t_rxd1[2][0] = 1350ns;
slave_timing[0][128+8].t_rxd2[0][2] = 1318ns;
slave_timing[0][128+8].t_rxd2[2][0] = 796ns;
slave_timing[0][128+8].t_rxd2[1][2] = 1047ns;
slave_timing[0][128+8].t_rxd2[2][1] = 1068ns;

slave_timing[0][128+9].info_corner          = 1;
slave_timing[0][128+9].info_temp__j__       = -40;
slave_timing[0][128+9].info_i__quite_rec__  = 0.003000000;
slave_timing[0][128+9].info_dtr__ib__       = -1;
slave_timing[0][128+9].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+9].info_i__max_slave__  = 0.025000000;
slave_timing[0][128+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][128+9].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+9].t_rxd1[0][1] = 1026ns;
slave_timing[0][128+9].t_rxd1[1][0] = 1112ns;
slave_timing[0][128+9].t_rxd1[0][2] = 768ns;
slave_timing[0][128+9].t_rxd1[2][0] = 1379ns;
slave_timing[0][128+9].t_rxd2[0][2] = 1224ns;
slave_timing[0][128+9].t_rxd2[2][0] = 848ns;
slave_timing[0][128+9].t_rxd2[1][2] = 928ns;
slave_timing[0][128+9].t_rxd2[2][1] = 1194ns;

slave_timing[0][128+10].info_corner          = 1;
slave_timing[0][128+10].info_temp__j__       = -40;
slave_timing[0][128+10].info_i__quite_rec__  = 0.003000000;
slave_timing[0][128+10].info_dtr__ib__       = 1;
slave_timing[0][128+10].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+10].info_i__max_slave__  = 0.023000000;
slave_timing[0][128+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][128+10].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+10].t_rxd1[0][1] = 1115ns;
slave_timing[0][128+10].t_rxd1[1][0] = 1042ns;
slave_timing[0][128+10].t_rxd1[0][2] = 814ns;
slave_timing[0][128+10].t_rxd1[2][0] = 1316ns;
slave_timing[0][128+10].t_rxd2[0][2] = 1430ns;
slave_timing[0][128+10].t_rxd2[2][0] = 738ns;
slave_timing[0][128+10].t_rxd2[1][2] = 1174ns;
slave_timing[0][128+10].t_rxd2[2][1] = 963ns;

slave_timing[0][128+11].info_corner          = 1;
slave_timing[0][128+11].info_temp__j__       = -40;
slave_timing[0][128+11].info_i__quite_rec__  = 0.003000000;
slave_timing[0][128+11].info_dtr__ib__       = 1;
slave_timing[0][128+11].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+11].info_i__max_slave__  = 0.025000000;
slave_timing[0][128+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][128+11].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+11].t_rxd1[0][1] = 1065ns;
slave_timing[0][128+11].t_rxd1[1][0] = 1077ns;
slave_timing[0][128+11].t_rxd1[0][2] = 790ns;
slave_timing[0][128+11].t_rxd1[2][0] = 1348ns;
slave_timing[0][128+11].t_rxd2[0][2] = 1305ns;
slave_timing[0][128+11].t_rxd2[2][0] = 802ns;
slave_timing[0][128+11].t_rxd2[1][2] = 1031ns;
slave_timing[0][128+11].t_rxd2[2][1] = 1080ns;

slave_timing[0][128+12].info_corner          = 1;
slave_timing[0][128+12].info_temp__j__       = -40;
slave_timing[0][128+12].info_i__quite_rec__  = 0.003000000;
slave_timing[0][128+12].info_dtr__ib__       = -1;
slave_timing[0][128+12].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+12].info_i__max_slave__  = 0.023000000;
slave_timing[0][128+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][128+12].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+12].t_rxd1[0][1] = 1152ns;
slave_timing[0][128+12].t_rxd1[1][0] = 1149ns;
slave_timing[0][128+12].t_rxd1[0][2] = 857ns;
slave_timing[0][128+12].t_rxd1[2][0] = 1415ns;
slave_timing[0][128+12].t_rxd2[0][2] = 1343ns;
slave_timing[0][128+12].t_rxd2[2][0] = 813ns;
slave_timing[0][128+12].t_rxd2[1][2] = 1058ns;
slave_timing[0][128+12].t_rxd2[2][1] = 1080ns;

slave_timing[0][128+13].info_corner          = 1;
slave_timing[0][128+13].info_temp__j__       = -40;
slave_timing[0][128+13].info_i__quite_rec__  = 0.003000000;
slave_timing[0][128+13].info_dtr__ib__       = -1;
slave_timing[0][128+13].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+13].info_i__max_slave__  = 0.025000000;
slave_timing[0][128+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][128+13].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+13].t_rxd1[0][1] = 1101ns;
slave_timing[0][128+13].t_rxd1[1][0] = 1183ns;
slave_timing[0][128+13].t_rxd1[0][2] = 832ns;
slave_timing[0][128+13].t_rxd1[2][0] = 1447ns;
slave_timing[0][128+13].t_rxd2[0][2] = 1249ns;
slave_timing[0][128+13].t_rxd2[2][0] = 869ns;
slave_timing[0][128+13].t_rxd2[1][2] = 940ns;
slave_timing[0][128+13].t_rxd2[2][1] = 1202ns;

slave_timing[0][128+14].info_corner          = 1;
slave_timing[0][128+14].info_temp__j__       = -40;
slave_timing[0][128+14].info_i__quite_rec__  = 0.003000000;
slave_timing[0][128+14].info_dtr__ib__       = 1;
slave_timing[0][128+14].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+14].info_i__max_slave__  = 0.023000000;
slave_timing[0][128+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][128+14].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+14].t_rxd1[0][1] = 1201ns;
slave_timing[0][128+14].t_rxd1[1][0] = 1111ns;
slave_timing[0][128+14].t_rxd1[0][2] = 877ns;
slave_timing[0][128+14].t_rxd1[2][0] = 1384ns;
slave_timing[0][128+14].t_rxd2[0][2] = 1451ns;
slave_timing[0][128+14].t_rxd2[2][0] = 760ns;
slave_timing[0][128+14].t_rxd2[1][2] = 1185ns;
slave_timing[0][128+14].t_rxd2[2][1] = 978ns;

slave_timing[0][128+15].info_corner          = 1;
slave_timing[0][128+15].info_temp__j__       = -40;
slave_timing[0][128+15].info_i__quite_rec__  = 0.003000000;
slave_timing[0][128+15].info_dtr__ib__       = 1;
slave_timing[0][128+15].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+15].info_i__max_slave__  = 0.025000000;
slave_timing[0][128+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][128+15].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+15].t_rxd1[0][1] = 1146ns;
slave_timing[0][128+15].t_rxd1[1][0] = 1150ns;
slave_timing[0][128+15].t_rxd1[0][2] = 853ns;
slave_timing[0][128+15].t_rxd1[2][0] = 1415ns;
slave_timing[0][128+15].t_rxd2[0][2] = 1328ns;
slave_timing[0][128+15].t_rxd2[2][0] = 821ns;
slave_timing[0][128+15].t_rxd2[1][2] = 1044ns;
slave_timing[0][128+15].t_rxd2[2][1] = 1095ns;

slave_timing[0][128+16].info_corner          = 1;
slave_timing[0][128+16].info_temp__j__       = -40;
slave_timing[0][128+16].info_i__quite_rec__  = 0.000000000;
slave_timing[0][128+16].info_dtr__ib__       = -1;
slave_timing[0][128+16].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+16].info_i__max_slave__  = 0.023000000;
slave_timing[0][128+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][128+16].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+16].t_rxd1[0][1] = 1063ns;
slave_timing[0][128+16].t_rxd1[1][0] = 1082ns;
slave_timing[0][128+16].t_rxd1[0][2] = 787ns;
slave_timing[0][128+16].t_rxd1[2][0] = 1352ns;
slave_timing[0][128+16].t_rxd2[0][2] = 1312ns;
slave_timing[0][128+16].t_rxd2[2][0] = 797ns;
slave_timing[0][128+16].t_rxd2[1][2] = 1043ns;
slave_timing[0][128+16].t_rxd2[2][1] = 1077ns;

slave_timing[0][128+17].info_corner          = 1;
slave_timing[0][128+17].info_temp__j__       = -40;
slave_timing[0][128+17].info_i__quite_rec__  = 0.000000000;
slave_timing[0][128+17].info_dtr__ib__       = -1;
slave_timing[0][128+17].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+17].info_i__max_slave__  = 0.025000000;
slave_timing[0][128+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][128+17].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+17].t_rxd1[0][1] = 1019ns;
slave_timing[0][128+17].t_rxd1[1][0] = 1117ns;
slave_timing[0][128+17].t_rxd1[0][2] = 764ns;
slave_timing[0][128+17].t_rxd1[2][0] = 1383ns;
slave_timing[0][128+17].t_rxd2[0][2] = 1219ns;
slave_timing[0][128+17].t_rxd2[2][0] = 850ns;
slave_timing[0][128+17].t_rxd2[1][2] = 924ns;
slave_timing[0][128+17].t_rxd2[2][1] = 1205ns;

slave_timing[0][128+18].info_corner          = 1;
slave_timing[0][128+18].info_temp__j__       = -40;
slave_timing[0][128+18].info_i__quite_rec__  = 0.000000000;
slave_timing[0][128+18].info_dtr__ib__       = 1;
slave_timing[0][128+18].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+18].info_i__max_slave__  = 0.023000000;
slave_timing[0][128+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][128+18].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+18].t_rxd1[0][1] = 1109ns;
slave_timing[0][128+18].t_rxd1[1][0] = 1048ns;
slave_timing[0][128+18].t_rxd1[0][2] = 808ns;
slave_timing[0][128+18].t_rxd1[2][0] = 1327ns;
slave_timing[0][128+18].t_rxd2[0][2] = 1417ns;
slave_timing[0][128+18].t_rxd2[2][0] = 744ns;
slave_timing[0][128+18].t_rxd2[1][2] = 1163ns;
slave_timing[0][128+18].t_rxd2[2][1] = 964ns;

slave_timing[0][128+19].info_corner          = 1;
slave_timing[0][128+19].info_temp__j__       = -40;
slave_timing[0][128+19].info_i__quite_rec__  = 0.000000000;
slave_timing[0][128+19].info_dtr__ib__       = 1;
slave_timing[0][128+19].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+19].info_i__max_slave__  = 0.025000000;
slave_timing[0][128+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][128+19].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+19].t_rxd1[0][1] = 1060ns;
slave_timing[0][128+19].t_rxd1[1][0] = 1088ns;
slave_timing[0][128+19].t_rxd1[0][2] = 787ns;
slave_timing[0][128+19].t_rxd1[2][0] = 1357ns;
slave_timing[0][128+19].t_rxd2[0][2] = 1297ns;
slave_timing[0][128+19].t_rxd2[2][0] = 802ns;
slave_timing[0][128+19].t_rxd2[1][2] = 1024ns;
slave_timing[0][128+19].t_rxd2[2][1] = 1085ns;

slave_timing[0][128+20].info_corner          = 1;
slave_timing[0][128+20].info_temp__j__       = -40;
slave_timing[0][128+20].info_i__quite_rec__  = 0.000000000;
slave_timing[0][128+20].info_dtr__ib__       = -1;
slave_timing[0][128+20].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+20].info_i__max_slave__  = 0.023000000;
slave_timing[0][128+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][128+20].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+20].t_rxd1[0][1] = 1145ns;
slave_timing[0][128+20].t_rxd1[1][0] = 1156ns;
slave_timing[0][128+20].t_rxd1[0][2] = 852ns;
slave_timing[0][128+20].t_rxd1[2][0] = 1421ns;
slave_timing[0][128+20].t_rxd2[0][2] = 1335ns;
slave_timing[0][128+20].t_rxd2[2][0] = 818ns;
slave_timing[0][128+20].t_rxd2[1][2] = 1053ns;
slave_timing[0][128+20].t_rxd2[2][1] = 1087ns;

slave_timing[0][128+21].info_corner          = 1;
slave_timing[0][128+21].info_temp__j__       = -40;
slave_timing[0][128+21].info_i__quite_rec__  = 0.000000000;
slave_timing[0][128+21].info_dtr__ib__       = -1;
slave_timing[0][128+21].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+21].info_i__max_slave__  = 0.025000000;
slave_timing[0][128+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][128+21].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+21].t_rxd1[0][1] = 1097ns;
slave_timing[0][128+21].t_rxd1[1][0] = 1189ns;
slave_timing[0][128+21].t_rxd1[0][2] = 828ns;
slave_timing[0][128+21].t_rxd1[2][0] = 1449ns;
slave_timing[0][128+21].t_rxd2[0][2] = 1244ns;
slave_timing[0][128+21].t_rxd2[2][0] = 869ns;
slave_timing[0][128+21].t_rxd2[1][2] = 935ns;
slave_timing[0][128+21].t_rxd2[2][1] = 1210ns;

slave_timing[0][128+22].info_corner          = 1;
slave_timing[0][128+22].info_temp__j__       = -40;
slave_timing[0][128+22].info_i__quite_rec__  = 0.000000000;
slave_timing[0][128+22].info_dtr__ib__       = 1;
slave_timing[0][128+22].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+22].info_i__max_slave__  = 0.023000000;
slave_timing[0][128+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][128+22].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+22].t_rxd1[0][1] = 1191ns;
slave_timing[0][128+22].t_rxd1[1][0] = 1123ns;
slave_timing[0][128+22].t_rxd1[0][2] = 874ns;
slave_timing[0][128+22].t_rxd1[2][0] = 1393ns;
slave_timing[0][128+22].t_rxd2[0][2] = 1439ns;
slave_timing[0][128+22].t_rxd2[2][0] = 759ns;
slave_timing[0][128+22].t_rxd2[1][2] = 1175ns;
slave_timing[0][128+22].t_rxd2[2][1] = 980ns;

slave_timing[0][128+23].info_corner          = 1;
slave_timing[0][128+23].info_temp__j__       = -40;
slave_timing[0][128+23].info_i__quite_rec__  = 0.000000000;
slave_timing[0][128+23].info_dtr__ib__       = 1;
slave_timing[0][128+23].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+23].info_i__max_slave__  = 0.025000000;
slave_timing[0][128+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][128+23].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+23].t_rxd1[0][1] = 1137ns;
slave_timing[0][128+23].t_rxd1[1][0] = 1159ns;
slave_timing[0][128+23].t_rxd1[0][2] = 848ns;
slave_timing[0][128+23].t_rxd1[2][0] = 1423ns;
slave_timing[0][128+23].t_rxd2[0][2] = 1318ns;
slave_timing[0][128+23].t_rxd2[2][0] = 820ns;
slave_timing[0][128+23].t_rxd2[1][2] = 1032ns;
slave_timing[0][128+23].t_rxd2[2][1] = 1097ns;

slave_timing[0][128+24].info_corner          = 1;
slave_timing[0][128+24].info_temp__j__       = -40;
slave_timing[0][128+24].info_i__quite_rec__  = 0.040000000;
slave_timing[0][128+24].info_dtr__ib__       = -1;
slave_timing[0][128+24].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+24].info_i__max_slave__  = 0.023000000;
slave_timing[0][128+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][128+24].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+24].t_rxd1[0][1] = 1067ns;
slave_timing[0][128+24].t_rxd1[1][0] = 1065ns;
slave_timing[0][128+24].t_rxd1[0][2] = 785ns;
slave_timing[0][128+24].t_rxd1[2][0] = 1334ns;
slave_timing[0][128+24].t_rxd2[0][2] = 1317ns;
slave_timing[0][128+24].t_rxd2[2][0] = 792ns;
slave_timing[0][128+24].t_rxd2[1][2] = 1053ns;
slave_timing[0][128+24].t_rxd2[2][1] = 1063ns;

slave_timing[0][128+25].info_corner          = 1;
slave_timing[0][128+25].info_temp__j__       = -40;
slave_timing[0][128+25].info_i__quite_rec__  = 0.040000000;
slave_timing[0][128+25].info_dtr__ib__       = -1;
slave_timing[0][128+25].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+25].info_i__max_slave__  = 0.025000000;
slave_timing[0][128+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][128+25].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+25].t_rxd1[0][1] = 1020ns;
slave_timing[0][128+25].t_rxd1[1][0] = 1096ns;
slave_timing[0][128+25].t_rxd1[0][2] = 763ns;
slave_timing[0][128+25].t_rxd1[2][0] = 1366ns;
slave_timing[0][128+25].t_rxd2[0][2] = 1224ns;
slave_timing[0][128+25].t_rxd2[2][0] = 847ns;
slave_timing[0][128+25].t_rxd2[1][2] = 930ns;
slave_timing[0][128+25].t_rxd2[2][1] = 1191ns;

slave_timing[0][128+26].info_corner          = 1;
slave_timing[0][128+26].info_temp__j__       = -40;
slave_timing[0][128+26].info_i__quite_rec__  = 0.040000000;
slave_timing[0][128+26].info_dtr__ib__       = 1;
slave_timing[0][128+26].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+26].info_i__max_slave__  = 0.023000000;
slave_timing[0][128+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][128+26].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+26].t_rxd1[0][1] = 1094ns;
slave_timing[0][128+26].t_rxd1[1][0] = 1043ns;
slave_timing[0][128+26].t_rxd1[0][2] = 801ns;
slave_timing[0][128+26].t_rxd1[2][0] = 1320ns;
slave_timing[0][128+26].t_rxd2[0][2] = 1415ns;
slave_timing[0][128+26].t_rxd2[2][0] = 749ns;
slave_timing[0][128+26].t_rxd2[1][2] = 1161ns;
slave_timing[0][128+26].t_rxd2[2][1] = 976ns;

slave_timing[0][128+27].info_corner          = 1;
slave_timing[0][128+27].info_temp__j__       = -40;
slave_timing[0][128+27].info_i__quite_rec__  = 0.040000000;
slave_timing[0][128+27].info_dtr__ib__       = 1;
slave_timing[0][128+27].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+27].info_i__max_slave__  = 0.025000000;
slave_timing[0][128+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][128+27].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+27].t_rxd1[0][1] = 1045ns;
slave_timing[0][128+27].t_rxd1[1][0] = 1080ns;
slave_timing[0][128+27].t_rxd1[0][2] = 777ns;
slave_timing[0][128+27].t_rxd1[2][0] = 1349ns;
slave_timing[0][128+27].t_rxd2[0][2] = 1293ns;
slave_timing[0][128+27].t_rxd2[2][0] = 805ns;
slave_timing[0][128+27].t_rxd2[1][2] = 1021ns;
slave_timing[0][128+27].t_rxd2[2][1] = 1094ns;

slave_timing[0][128+28].info_corner          = 1;
slave_timing[0][128+28].info_temp__j__       = -40;
slave_timing[0][128+28].info_i__quite_rec__  = 0.040000000;
slave_timing[0][128+28].info_dtr__ib__       = -1;
slave_timing[0][128+28].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+28].info_i__max_slave__  = 0.023000000;
slave_timing[0][128+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][128+28].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+28].t_rxd1[0][1] = 1108ns;
slave_timing[0][128+28].t_rxd1[1][0] = 1109ns;
slave_timing[0][128+28].t_rxd1[0][2] = 824ns;
slave_timing[0][128+28].t_rxd1[2][0] = 1373ns;
slave_timing[0][128+28].t_rxd2[0][2] = 1331ns;
slave_timing[0][128+28].t_rxd2[2][0] = 810ns;
slave_timing[0][128+28].t_rxd2[1][2] = 1061ns;
slave_timing[0][128+28].t_rxd2[2][1] = 1078ns;

slave_timing[0][128+29].info_corner          = 1;
slave_timing[0][128+29].info_temp__j__       = -40;
slave_timing[0][128+29].info_i__quite_rec__  = 0.040000000;
slave_timing[0][128+29].info_dtr__ib__       = -1;
slave_timing[0][128+29].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+29].info_i__max_slave__  = 0.025000000;
slave_timing[0][128+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][128+29].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+29].t_rxd1[0][1] = 1062ns;
slave_timing[0][128+29].t_rxd1[1][0] = 1142ns;
slave_timing[0][128+29].t_rxd1[0][2] = 800ns;
slave_timing[0][128+29].t_rxd1[2][0] = 1401ns;
slave_timing[0][128+29].t_rxd2[0][2] = 1236ns;
slave_timing[0][128+29].t_rxd2[2][0] = 863ns;
slave_timing[0][128+29].t_rxd2[1][2] = 945ns;
slave_timing[0][128+29].t_rxd2[2][1] = 1199ns;

slave_timing[0][128+30].info_corner          = 1;
slave_timing[0][128+30].info_temp__j__       = -40;
slave_timing[0][128+30].info_i__quite_rec__  = 0.040000000;
slave_timing[0][128+30].info_dtr__ib__       = 1;
slave_timing[0][128+30].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+30].info_i__max_slave__  = 0.023000000;
slave_timing[0][128+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][128+30].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+30].t_rxd1[0][1] = 1141ns;
slave_timing[0][128+30].t_rxd1[1][0] = 1092ns;
slave_timing[0][128+30].t_rxd1[0][2] = 842ns;
slave_timing[0][128+30].t_rxd1[2][0] = 1358ns;
slave_timing[0][128+30].t_rxd2[0][2] = 1428ns;
slave_timing[0][128+30].t_rxd2[2][0] = 766ns;
slave_timing[0][128+30].t_rxd2[1][2] = 1171ns;
slave_timing[0][128+30].t_rxd2[2][1] = 989ns;

slave_timing[0][128+31].info_corner          = 1;
slave_timing[0][128+31].info_temp__j__       = -40;
slave_timing[0][128+31].info_i__quite_rec__  = 0.040000000;
slave_timing[0][128+31].info_dtr__ib__       = 1;
slave_timing[0][128+31].info_i__offset_rec__ = 0.000000000;
slave_timing[0][128+31].info_i__max_slave__  = 0.025000000;
slave_timing[0][128+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][128+31].info_r__dsi_bus__    = 5.000;

slave_timing[0][128+31].t_rxd1[0][1] = 1090ns;
slave_timing[0][128+31].t_rxd1[1][0] = 1126ns;
slave_timing[0][128+31].t_rxd1[0][2] = 817ns;
slave_timing[0][128+31].t_rxd1[2][0] = 1386ns;
slave_timing[0][128+31].t_rxd2[0][2] = 1307ns;
slave_timing[0][128+31].t_rxd2[2][0] = 821ns;
slave_timing[0][128+31].t_rxd2[1][2] = 1030ns;
slave_timing[0][128+31].t_rxd2[2][1] = 1098ns;

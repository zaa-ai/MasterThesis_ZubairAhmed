
`timescale 1ns/1ns

module pure_delay #(
    parameter DOMAIN_3V0 = 0
  )(
    input  i_a,
    output o_y
  );

  BUFFD1BWP7T delay_inst(
    .I (i_a),
    .Z (o_y)
  );

endmodule


import addresses_pkg::*;
import test_addresses_pkg::*;
import edf_epm_model_pkg::*;
import M52144A_pattern_pkg::*;
import ECC_pkg::*;

`include "dsi3_transaction_recorder.svh"
`include "dsi3_master_configuration_listener.svh"
`include "register_resetter.svh"
`include "chip_time_iterator.svh"

virtual clk_reset_if vif_clk_rst;

pdcm_buffer_writer_action_e action;

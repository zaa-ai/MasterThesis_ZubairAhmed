//-----------------------------------------------------------------------------
// Copyright (c) 2023 Elmos SE
// Author     : Eugene - Easy UVM Generator
//
// Description: This file has been generated automatically by Eugene
//				This file should not be modified manually. 
//-----------------------------------------------------------------------------
`ifndef REAL_SIGNAL_CONFIG_SV
`define REAL_SIGNAL_CONFIG_SV

// You can insert code here by setting agent_config_inc_before_class in file real_signal.tpl

class real_signal_config extends uvm_object;

	// Do not register config class with the factory
	
	virtual	real_signal_if vif;
	
	uvm_active_passive_enum is_active = UVM_ACTIVE;
	bit	coverage_enable;       
	
	real init_value = 0.0;
	time time_scale = 1ns;
	real value_scale = 0.01;
	
	// You can remove new by setting agent_config_generate_methods_inside_class = no in file real_signal.tpl
	function new(string name = "");
		super.new("real_signal_config");
	endfunction
	
	// You can insert code here by setting agent_config_inc_inside_class in file real_signal.tpl

endclass 

// You can insert code here by setting agent_config_inc_after_class in file real_signal.tpl

`endif

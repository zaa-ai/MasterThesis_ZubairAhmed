
slave_timing[2][32+0].info_corner          = 2;
slave_timing[2][32+0].info_temp__j__       = 125;
slave_timing[2][32+0].info_i__quite_rec__  = 0.006000000;
slave_timing[2][32+0].info_dtr__ib__       = -1;
slave_timing[2][32+0].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+0].info_i__max_slave__  = 0.023000000;
slave_timing[2][32+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][32+0].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+0].t_rxd1[0][1] = 2209ns;
slave_timing[2][32+0].t_rxd1[1][0] = 2237ns;
slave_timing[2][32+0].t_rxd1[0][2] = 1673ns;
slave_timing[2][32+0].t_rxd1[2][0] = 2700ns;
slave_timing[2][32+0].t_rxd2[0][2] = 2650ns;
slave_timing[2][32+0].t_rxd2[2][0] = 1684ns;
slave_timing[2][32+0].t_rxd2[1][2] = 2202ns;
slave_timing[2][32+0].t_rxd2[2][1] = 2213ns;

slave_timing[2][32+1].info_corner          = 2;
slave_timing[2][32+1].info_temp__j__       = 125;
slave_timing[2][32+1].info_i__quite_rec__  = 0.006000000;
slave_timing[2][32+1].info_dtr__ib__       = -1;
slave_timing[2][32+1].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+1].info_i__max_slave__  = 0.025000000;
slave_timing[2][32+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][32+1].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+1].t_rxd1[0][1] = 2114ns;
slave_timing[2][32+1].t_rxd1[1][0] = 2301ns;
slave_timing[2][32+1].t_rxd1[0][2] = 1621ns;
slave_timing[2][32+1].t_rxd1[2][0] = 2740ns;
slave_timing[2][32+1].t_rxd2[0][2] = 2499ns;
slave_timing[2][32+1].t_rxd2[2][0] = 1799ns;
slave_timing[2][32+1].t_rxd2[1][2] = 1976ns;
slave_timing[2][32+1].t_rxd2[2][1] = 2438ns;

slave_timing[2][32+2].info_corner          = 2;
slave_timing[2][32+2].info_temp__j__       = 125;
slave_timing[2][32+2].info_i__quite_rec__  = 0.006000000;
slave_timing[2][32+2].info_dtr__ib__       = 1;
slave_timing[2][32+2].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+2].info_i__max_slave__  = 0.023000000;
slave_timing[2][32+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][32+2].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+2].t_rxd1[0][1] = 2249ns;
slave_timing[2][32+2].t_rxd1[1][0] = 2173ns;
slave_timing[2][32+2].t_rxd1[0][2] = 1694ns;
slave_timing[2][32+2].t_rxd1[2][0] = 2651ns;
slave_timing[2][32+2].t_rxd2[0][2] = 2780ns;
slave_timing[2][32+2].t_rxd2[2][0] = 1576ns;
slave_timing[2][32+2].t_rxd2[1][2] = 2388ns;
slave_timing[2][32+2].t_rxd2[2][1] = 2029ns;

slave_timing[2][32+3].info_corner          = 2;
slave_timing[2][32+3].info_temp__j__       = 125;
slave_timing[2][32+3].info_i__quite_rec__  = 0.006000000;
slave_timing[2][32+3].info_dtr__ib__       = 1;
slave_timing[2][32+3].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+3].info_i__max_slave__  = 0.025000000;
slave_timing[2][32+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][32+3].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+3].t_rxd1[0][1] = 2167ns;
slave_timing[2][32+3].t_rxd1[1][0] = 2246ns;
slave_timing[2][32+3].t_rxd1[0][2] = 1644ns;
slave_timing[2][32+3].t_rxd1[2][0] = 2693ns;
slave_timing[2][32+3].t_rxd2[0][2] = 2600ns;
slave_timing[2][32+3].t_rxd2[2][0] = 1706ns;
slave_timing[2][32+3].t_rxd2[1][2] = 2129ns;
slave_timing[2][32+3].t_rxd2[2][1] = 2253ns;

slave_timing[2][32+4].info_corner          = 2;
slave_timing[2][32+4].info_temp__j__       = 125;
slave_timing[2][32+4].info_i__quite_rec__  = 0.006000000;
slave_timing[2][32+4].info_dtr__ib__       = -1;
slave_timing[2][32+4].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+4].info_i__max_slave__  = 0.023000000;
slave_timing[2][32+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][32+4].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+4].t_rxd1[0][1] = 2370ns;
slave_timing[2][32+4].t_rxd1[1][0] = 2361ns;
slave_timing[2][32+4].t_rxd1[0][2] = 1793ns;
slave_timing[2][32+4].t_rxd1[2][0] = 2829ns;
slave_timing[2][32+4].t_rxd2[0][2] = 2655ns;
slave_timing[2][32+4].t_rxd2[2][0] = 1712ns;
slave_timing[2][32+4].t_rxd2[1][2] = 2223ns;
slave_timing[2][32+4].t_rxd2[2][1] = 2237ns;

slave_timing[2][32+5].info_corner          = 2;
slave_timing[2][32+5].info_temp__j__       = 125;
slave_timing[2][32+5].info_i__quite_rec__  = 0.006000000;
slave_timing[2][32+5].info_dtr__ib__       = -1;
slave_timing[2][32+5].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+5].info_i__max_slave__  = 0.025000000;
slave_timing[2][32+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][32+5].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+5].t_rxd1[0][1] = 2282ns;
slave_timing[2][32+5].t_rxd1[1][0] = 2437ns;
slave_timing[2][32+5].t_rxd1[0][2] = 1763ns;
slave_timing[2][32+5].t_rxd1[2][0] = 2864ns;
slave_timing[2][32+5].t_rxd2[0][2] = 2533ns;
slave_timing[2][32+5].t_rxd2[2][0] = 1825ns;
slave_timing[2][32+5].t_rxd2[1][2] = 1998ns;
slave_timing[2][32+5].t_rxd2[2][1] = 2431ns;

slave_timing[2][32+6].info_corner          = 2;
slave_timing[2][32+6].info_temp__j__       = 125;
slave_timing[2][32+6].info_i__quite_rec__  = 0.006000000;
slave_timing[2][32+6].info_dtr__ib__       = 1;
slave_timing[2][32+6].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+6].info_i__max_slave__  = 0.023000000;
slave_timing[2][32+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][32+6].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+6].t_rxd1[0][1] = 2416ns;
slave_timing[2][32+6].t_rxd1[1][0] = 2316ns;
slave_timing[2][32+6].t_rxd1[0][2] = 1836ns;
slave_timing[2][32+6].t_rxd1[2][0] = 2777ns;
slave_timing[2][32+6].t_rxd2[0][2] = 2806ns;
slave_timing[2][32+6].t_rxd2[2][0] = 1603ns;
slave_timing[2][32+6].t_rxd2[1][2] = 2404ns;
slave_timing[2][32+6].t_rxd2[2][1] = 2057ns;

slave_timing[2][32+7].info_corner          = 2;
slave_timing[2][32+7].info_temp__j__       = 125;
slave_timing[2][32+7].info_i__quite_rec__  = 0.006000000;
slave_timing[2][32+7].info_dtr__ib__       = 1;
slave_timing[2][32+7].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+7].info_i__max_slave__  = 0.025000000;
slave_timing[2][32+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][32+7].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+7].t_rxd1[0][1] = 2322ns;
slave_timing[2][32+7].t_rxd1[1][0] = 2377ns;
slave_timing[2][32+7].t_rxd1[0][2] = 1782ns;
slave_timing[2][32+7].t_rxd1[2][0] = 2822ns;
slave_timing[2][32+7].t_rxd2[0][2] = 2631ns;
slave_timing[2][32+7].t_rxd2[2][0] = 1734ns;
slave_timing[2][32+7].t_rxd2[1][2] = 2152ns;
slave_timing[2][32+7].t_rxd2[2][1] = 2250ns;

slave_timing[2][32+8].info_corner          = 2;
slave_timing[2][32+8].info_temp__j__       = 125;
slave_timing[2][32+8].info_i__quite_rec__  = 0.003000000;
slave_timing[2][32+8].info_dtr__ib__       = -1;
slave_timing[2][32+8].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+8].info_i__max_slave__  = 0.023000000;
slave_timing[2][32+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][32+8].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+8].t_rxd1[0][1] = 2190ns;
slave_timing[2][32+8].t_rxd1[1][0] = 2208ns;
slave_timing[2][32+8].t_rxd1[0][2] = 1658ns;
slave_timing[2][32+8].t_rxd1[2][0] = 2668ns;
slave_timing[2][32+8].t_rxd2[0][2] = 2647ns;
slave_timing[2][32+8].t_rxd2[2][0] = 1664ns;
slave_timing[2][32+8].t_rxd2[1][2] = 2204ns;
slave_timing[2][32+8].t_rxd2[2][1] = 2156ns;

slave_timing[2][32+9].info_corner          = 2;
slave_timing[2][32+9].info_temp__j__       = 125;
slave_timing[2][32+9].info_i__quite_rec__  = 0.003000000;
slave_timing[2][32+9].info_dtr__ib__       = -1;
slave_timing[2][32+9].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+9].info_i__max_slave__  = 0.025000000;
slave_timing[2][32+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][32+9].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+9].t_rxd1[0][1] = 2110ns;
slave_timing[2][32+9].t_rxd1[1][0] = 2267ns;
slave_timing[2][32+9].t_rxd1[0][2] = 1613ns;
slave_timing[2][32+9].t_rxd1[2][0] = 2711ns;
slave_timing[2][32+9].t_rxd2[0][2] = 2497ns;
slave_timing[2][32+9].t_rxd2[2][0] = 1780ns;
slave_timing[2][32+9].t_rxd2[1][2] = 1972ns;
slave_timing[2][32+9].t_rxd2[2][1] = 2415ns;

slave_timing[2][32+10].info_corner          = 2;
slave_timing[2][32+10].info_temp__j__       = 125;
slave_timing[2][32+10].info_i__quite_rec__  = 0.003000000;
slave_timing[2][32+10].info_dtr__ib__       = 1;
slave_timing[2][32+10].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+10].info_i__max_slave__  = 0.023000000;
slave_timing[2][32+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][32+10].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+10].t_rxd1[0][1] = 2232ns;
slave_timing[2][32+10].t_rxd1[1][0] = 2114ns;
slave_timing[2][32+10].t_rxd1[0][2] = 1676ns;
slave_timing[2][32+10].t_rxd1[2][0] = 2604ns;
slave_timing[2][32+10].t_rxd2[0][2] = 2770ns;
slave_timing[2][32+10].t_rxd2[2][0] = 1559ns;
slave_timing[2][32+10].t_rxd2[1][2] = 2394ns;
slave_timing[2][32+10].t_rxd2[2][1] = 2007ns;

slave_timing[2][32+11].info_corner          = 2;
slave_timing[2][32+11].info_temp__j__       = 125;
slave_timing[2][32+11].info_i__quite_rec__  = 0.003000000;
slave_timing[2][32+11].info_dtr__ib__       = 1;
slave_timing[2][32+11].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+11].info_i__max_slave__  = 0.025000000;
slave_timing[2][32+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][32+11].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+11].t_rxd1[0][1] = 2149ns;
slave_timing[2][32+11].t_rxd1[1][0] = 2200ns;
slave_timing[2][32+11].t_rxd1[0][2] = 1623ns;
slave_timing[2][32+11].t_rxd1[2][0] = 2649ns;
slave_timing[2][32+11].t_rxd2[0][2] = 2586ns;
slave_timing[2][32+11].t_rxd2[2][0] = 1687ns;
slave_timing[2][32+11].t_rxd2[1][2] = 2129ns;
slave_timing[2][32+11].t_rxd2[2][1] = 2233ns;

slave_timing[2][32+12].info_corner          = 2;
slave_timing[2][32+12].info_temp__j__       = 125;
slave_timing[2][32+12].info_i__quite_rec__  = 0.003000000;
slave_timing[2][32+12].info_dtr__ib__       = -1;
slave_timing[2][32+12].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+12].info_i__max_slave__  = 0.023000000;
slave_timing[2][32+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][32+12].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+12].t_rxd1[0][1] = 2366ns;
slave_timing[2][32+12].t_rxd1[1][0] = 2339ns;
slave_timing[2][32+12].t_rxd1[0][2] = 1810ns;
slave_timing[2][32+12].t_rxd1[2][0] = 2794ns;
slave_timing[2][32+12].t_rxd2[0][2] = 2677ns;
slave_timing[2][32+12].t_rxd2[2][0] = 1694ns;
slave_timing[2][32+12].t_rxd2[1][2] = 2224ns;
slave_timing[2][32+12].t_rxd2[2][1] = 2198ns;

slave_timing[2][32+13].info_corner          = 2;
slave_timing[2][32+13].info_temp__j__       = 125;
slave_timing[2][32+13].info_i__quite_rec__  = 0.003000000;
slave_timing[2][32+13].info_dtr__ib__       = -1;
slave_timing[2][32+13].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+13].info_i__max_slave__  = 0.025000000;
slave_timing[2][32+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][32+13].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+13].t_rxd1[0][1] = 2284ns;
slave_timing[2][32+13].t_rxd1[1][0] = 2408ns;
slave_timing[2][32+13].t_rxd1[0][2] = 1742ns;
slave_timing[2][32+13].t_rxd1[2][0] = 2838ns;
slave_timing[2][32+13].t_rxd2[0][2] = 2502ns;
slave_timing[2][32+13].t_rxd2[2][0] = 1807ns;
slave_timing[2][32+13].t_rxd2[1][2] = 1996ns;
slave_timing[2][32+13].t_rxd2[2][1] = 2432ns;

slave_timing[2][32+14].info_corner          = 2;
slave_timing[2][32+14].info_temp__j__       = 125;
slave_timing[2][32+14].info_i__quite_rec__  = 0.003000000;
slave_timing[2][32+14].info_dtr__ib__       = 1;
slave_timing[2][32+14].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+14].info_i__max_slave__  = 0.023000000;
slave_timing[2][32+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][32+14].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+14].t_rxd1[0][1] = 2414ns;
slave_timing[2][32+14].t_rxd1[1][0] = 2266ns;
slave_timing[2][32+14].t_rxd1[0][2] = 1828ns;
slave_timing[2][32+14].t_rxd1[2][0] = 2730ns;
slave_timing[2][32+14].t_rxd2[0][2] = 2794ns;
slave_timing[2][32+14].t_rxd2[2][0] = 1586ns;
slave_timing[2][32+14].t_rxd2[1][2] = 2407ns;
slave_timing[2][32+14].t_rxd2[2][1] = 2020ns;

slave_timing[2][32+15].info_corner          = 2;
slave_timing[2][32+15].info_temp__j__       = 125;
slave_timing[2][32+15].info_i__quite_rec__  = 0.003000000;
slave_timing[2][32+15].info_dtr__ib__       = 1;
slave_timing[2][32+15].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+15].info_i__max_slave__  = 0.025000000;
slave_timing[2][32+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][32+15].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+15].t_rxd1[0][1] = 2318ns;
slave_timing[2][32+15].t_rxd1[1][0] = 2331ns;
slave_timing[2][32+15].t_rxd1[0][2] = 1777ns;
slave_timing[2][32+15].t_rxd1[2][0] = 2771ns;
slave_timing[2][32+15].t_rxd2[0][2] = 2615ns;
slave_timing[2][32+15].t_rxd2[2][0] = 1716ns;
slave_timing[2][32+15].t_rxd2[1][2] = 2154ns;
slave_timing[2][32+15].t_rxd2[2][1] = 2253ns;

slave_timing[2][32+16].info_corner          = 2;
slave_timing[2][32+16].info_temp__j__       = 125;
slave_timing[2][32+16].info_i__quite_rec__  = 0.000000000;
slave_timing[2][32+16].info_dtr__ib__       = -1;
slave_timing[2][32+16].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+16].info_i__max_slave__  = 0.023000000;
slave_timing[2][32+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][32+16].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+16].t_rxd1[0][1] = 2176ns;
slave_timing[2][32+16].t_rxd1[1][0] = 2154ns;
slave_timing[2][32+16].t_rxd1[0][2] = 1636ns;
slave_timing[2][32+16].t_rxd1[2][0] = 2621ns;
slave_timing[2][32+16].t_rxd2[0][2] = 2630ns;
slave_timing[2][32+16].t_rxd2[2][0] = 1647ns;
slave_timing[2][32+16].t_rxd2[1][2] = 2199ns;
slave_timing[2][32+16].t_rxd2[2][1] = 2156ns;

slave_timing[2][32+17].info_corner          = 2;
slave_timing[2][32+17].info_temp__j__       = 125;
slave_timing[2][32+17].info_i__quite_rec__  = 0.000000000;
slave_timing[2][32+17].info_dtr__ib__       = -1;
slave_timing[2][32+17].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+17].info_i__max_slave__  = 0.025000000;
slave_timing[2][32+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][32+17].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+17].t_rxd1[0][1] = 2091ns;
slave_timing[2][32+17].t_rxd1[1][0] = 2221ns;
slave_timing[2][32+17].t_rxd1[0][2] = 1592ns;
slave_timing[2][32+17].t_rxd1[2][0] = 2663ns;
slave_timing[2][32+17].t_rxd2[0][2] = 2474ns;
slave_timing[2][32+17].t_rxd2[2][0] = 1763ns;
slave_timing[2][32+17].t_rxd2[1][2] = 1976ns;
slave_timing[2][32+17].t_rxd2[2][1] = 2387ns;

slave_timing[2][32+18].info_corner          = 2;
slave_timing[2][32+18].info_temp__j__       = 125;
slave_timing[2][32+18].info_i__quite_rec__  = 0.000000000;
slave_timing[2][32+18].info_dtr__ib__       = 1;
slave_timing[2][32+18].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+18].info_i__max_slave__  = 0.023000000;
slave_timing[2][32+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][32+18].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+18].t_rxd1[0][1] = 2215ns;
slave_timing[2][32+18].t_rxd1[1][0] = 2094ns;
slave_timing[2][32+18].t_rxd1[0][2] = 1656ns;
slave_timing[2][32+18].t_rxd1[2][0] = 2567ns;
slave_timing[2][32+18].t_rxd2[0][2] = 2747ns;
slave_timing[2][32+18].t_rxd2[2][0] = 1532ns;
slave_timing[2][32+18].t_rxd2[1][2] = 2381ns;
slave_timing[2][32+18].t_rxd2[2][1] = 1933ns;

slave_timing[2][32+19].info_corner          = 2;
slave_timing[2][32+19].info_temp__j__       = 125;
slave_timing[2][32+19].info_i__quite_rec__  = 0.000000000;
slave_timing[2][32+19].info_dtr__ib__       = 1;
slave_timing[2][32+19].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+19].info_i__max_slave__  = 0.025000000;
slave_timing[2][32+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][32+19].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+19].t_rxd1[0][1] = 2131ns;
slave_timing[2][32+19].t_rxd1[1][0] = 2172ns;
slave_timing[2][32+19].t_rxd1[0][2] = 1607ns;
slave_timing[2][32+19].t_rxd1[2][0] = 2611ns;
slave_timing[2][32+19].t_rxd2[0][2] = 2560ns;
slave_timing[2][32+19].t_rxd2[2][0] = 1663ns;
slave_timing[2][32+19].t_rxd2[1][2] = 2118ns;
slave_timing[2][32+19].t_rxd2[2][1] = 2191ns;

slave_timing[2][32+20].info_corner          = 2;
slave_timing[2][32+20].info_temp__j__       = 125;
slave_timing[2][32+20].info_i__quite_rec__  = 0.000000000;
slave_timing[2][32+20].info_dtr__ib__       = -1;
slave_timing[2][32+20].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+20].info_i__max_slave__  = 0.023000000;
slave_timing[2][32+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][32+20].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+20].t_rxd1[0][1] = 2356ns;
slave_timing[2][32+20].t_rxd1[1][0] = 2298ns;
slave_timing[2][32+20].t_rxd1[0][2] = 1804ns;
slave_timing[2][32+20].t_rxd1[2][0] = 2743ns;
slave_timing[2][32+20].t_rxd2[0][2] = 2653ns;
slave_timing[2][32+20].t_rxd2[2][0] = 1671ns;
slave_timing[2][32+20].t_rxd2[1][2] = 2214ns;
slave_timing[2][32+20].t_rxd2[2][1] = 2161ns;

slave_timing[2][32+21].info_corner          = 2;
slave_timing[2][32+21].info_temp__j__       = 125;
slave_timing[2][32+21].info_i__quite_rec__  = 0.000000000;
slave_timing[2][32+21].info_dtr__ib__       = -1;
slave_timing[2][32+21].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+21].info_i__max_slave__  = 0.025000000;
slave_timing[2][32+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][32+21].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+21].t_rxd1[0][1] = 2273ns;
slave_timing[2][32+21].t_rxd1[1][0] = 2360ns;
slave_timing[2][32+21].t_rxd1[0][2] = 1754ns;
slave_timing[2][32+21].t_rxd1[2][0] = 2786ns;
slave_timing[2][32+21].t_rxd2[0][2] = 2501ns;
slave_timing[2][32+21].t_rxd2[2][0] = 1788ns;
slave_timing[2][32+21].t_rxd2[1][2] = 2031ns;
slave_timing[2][32+21].t_rxd2[2][1] = 2373ns;

slave_timing[2][32+22].info_corner          = 2;
slave_timing[2][32+22].info_temp__j__       = 125;
slave_timing[2][32+22].info_i__quite_rec__  = 0.000000000;
slave_timing[2][32+22].info_dtr__ib__       = 1;
slave_timing[2][32+22].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+22].info_i__max_slave__  = 0.023000000;
slave_timing[2][32+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][32+22].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+22].t_rxd1[0][1] = 2402ns;
slave_timing[2][32+22].t_rxd1[1][0] = 2237ns;
slave_timing[2][32+22].t_rxd1[0][2] = 1822ns;
slave_timing[2][32+22].t_rxd1[2][0] = 2696ns;
slave_timing[2][32+22].t_rxd2[0][2] = 2764ns;
slave_timing[2][32+22].t_rxd2[2][0] = 1530ns;
slave_timing[2][32+22].t_rxd2[1][2] = 2432ns;
slave_timing[2][32+22].t_rxd2[2][1] = 1936ns;

slave_timing[2][32+23].info_corner          = 2;
slave_timing[2][32+23].info_temp__j__       = 125;
slave_timing[2][32+23].info_i__quite_rec__  = 0.000000000;
slave_timing[2][32+23].info_dtr__ib__       = 1;
slave_timing[2][32+23].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+23].info_i__max_slave__  = 0.025000000;
slave_timing[2][32+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][32+23].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+23].t_rxd1[0][1] = 2309ns;
slave_timing[2][32+23].t_rxd1[1][0] = 2302ns;
slave_timing[2][32+23].t_rxd1[0][2] = 1772ns;
slave_timing[2][32+23].t_rxd1[2][0] = 2734ns;
slave_timing[2][32+23].t_rxd2[0][2] = 2586ns;
slave_timing[2][32+23].t_rxd2[2][0] = 1687ns;
slave_timing[2][32+23].t_rxd2[1][2] = 2138ns;
slave_timing[2][32+23].t_rxd2[2][1] = 2187ns;

slave_timing[2][32+24].info_corner          = 2;
slave_timing[2][32+24].info_temp__j__       = 125;
slave_timing[2][32+24].info_i__quite_rec__  = 0.040000000;
slave_timing[2][32+24].info_dtr__ib__       = -1;
slave_timing[2][32+24].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+24].info_i__max_slave__  = 0.023000000;
slave_timing[2][32+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][32+24].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+24].t_rxd1[0][1] = 2189ns;
slave_timing[2][32+24].t_rxd1[1][0] = 2245ns;
slave_timing[2][32+24].t_rxd1[0][2] = 1670ns;
slave_timing[2][32+24].t_rxd1[2][0] = 2702ns;
slave_timing[2][32+24].t_rxd2[0][2] = 2836ns;
slave_timing[2][32+24].t_rxd2[2][0] = 1849ns;
slave_timing[2][32+24].t_rxd2[1][2] = 2391ns;
slave_timing[2][32+24].t_rxd2[2][1] = 2413ns;

slave_timing[2][32+25].info_corner          = 2;
slave_timing[2][32+25].info_temp__j__       = 125;
slave_timing[2][32+25].info_i__quite_rec__  = 0.040000000;
slave_timing[2][32+25].info_dtr__ib__       = -1;
slave_timing[2][32+25].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+25].info_i__max_slave__  = 0.025000000;
slave_timing[2][32+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][32+25].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+25].t_rxd1[0][1] = 2109ns;
slave_timing[2][32+25].t_rxd1[1][0] = 2307ns;
slave_timing[2][32+25].t_rxd1[0][2] = 1622ns;
slave_timing[2][32+25].t_rxd1[2][0] = 2741ns;
slave_timing[2][32+25].t_rxd2[0][2] = 2677ns;
slave_timing[2][32+25].t_rxd2[2][0] = 1964ns;
slave_timing[2][32+25].t_rxd2[1][2] = 2181ns;
slave_timing[2][32+25].t_rxd2[2][1] = 2614ns;

slave_timing[2][32+26].info_corner          = 2;
slave_timing[2][32+26].info_temp__j__       = 125;
slave_timing[2][32+26].info_i__quite_rec__  = 0.040000000;
slave_timing[2][32+26].info_dtr__ib__       = 1;
slave_timing[2][32+26].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+26].info_i__max_slave__  = 0.023000000;
slave_timing[2][32+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][32+26].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+26].t_rxd1[0][1] = 2278ns;
slave_timing[2][32+26].t_rxd1[1][0] = 2160ns;
slave_timing[2][32+26].t_rxd1[0][2] = 1715ns;
slave_timing[2][32+26].t_rxd1[2][0] = 2645ns;
slave_timing[2][32+26].t_rxd2[0][2] = 2989ns;
slave_timing[2][32+26].t_rxd2[2][0] = 1730ns;
slave_timing[2][32+26].t_rxd2[1][2] = 2611ns;
slave_timing[2][32+26].t_rxd2[2][1] = 2196ns;

slave_timing[2][32+27].info_corner          = 2;
slave_timing[2][32+27].info_temp__j__       = 125;
slave_timing[2][32+27].info_i__quite_rec__  = 0.040000000;
slave_timing[2][32+27].info_dtr__ib__       = 1;
slave_timing[2][32+27].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+27].info_i__max_slave__  = 0.025000000;
slave_timing[2][32+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][32+27].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+27].t_rxd1[0][1] = 2198ns;
slave_timing[2][32+27].t_rxd1[1][0] = 2239ns;
slave_timing[2][32+27].t_rxd1[0][2] = 1665ns;
slave_timing[2][32+27].t_rxd1[2][0] = 2694ns;
slave_timing[2][32+27].t_rxd2[0][2] = 2802ns;
slave_timing[2][32+27].t_rxd2[2][0] = 1864ns;
slave_timing[2][32+27].t_rxd2[1][2] = 2346ns;
slave_timing[2][32+27].t_rxd2[2][1] = 2445ns;

slave_timing[2][32+28].info_corner          = 2;
slave_timing[2][32+28].info_temp__j__       = 125;
slave_timing[2][32+28].info_i__quite_rec__  = 0.040000000;
slave_timing[2][32+28].info_dtr__ib__       = -1;
slave_timing[2][32+28].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+28].info_i__max_slave__  = 0.023000000;
slave_timing[2][32+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][32+28].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+28].t_rxd1[0][1] = 2257ns;
slave_timing[2][32+28].t_rxd1[1][0] = 2289ns;
slave_timing[2][32+28].t_rxd1[0][2] = 1723ns;
slave_timing[2][32+28].t_rxd1[2][0] = 2968ns;
slave_timing[2][32+28].t_rxd2[0][2] = 3314ns;
slave_timing[2][32+28].t_rxd2[2][0] = 2378ns;
slave_timing[2][32+28].t_rxd2[1][2] = 2969ns;
slave_timing[2][32+28].t_rxd2[2][1] = 3170ns;

slave_timing[2][32+29].info_corner          = 2;
slave_timing[2][32+29].info_temp__j__       = 125;
slave_timing[2][32+29].info_i__quite_rec__  = 0.040000000;
slave_timing[2][32+29].info_dtr__ib__       = -1;
slave_timing[2][32+29].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+29].info_i__max_slave__  = 0.025000000;
slave_timing[2][32+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][32+29].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+29].t_rxd1[0][1] = 2189ns;
slave_timing[2][32+29].t_rxd1[1][0] = 2359ns;
slave_timing[2][32+29].t_rxd1[0][2] = 1696ns;
slave_timing[2][32+29].t_rxd1[2][0] = 3079ns;
slave_timing[2][32+29].t_rxd2[0][2] = 3145ns;
slave_timing[2][32+29].t_rxd2[2][0] = 2539ns;
slave_timing[2][32+29].t_rxd2[1][2] = 2684ns;
slave_timing[2][32+29].t_rxd2[2][1] = 3515ns;

slave_timing[2][32+30].info_corner          = 2;
slave_timing[2][32+30].info_temp__j__       = 125;
slave_timing[2][32+30].info_i__quite_rec__  = 0.040000000;
slave_timing[2][32+30].info_dtr__ib__       = 1;
slave_timing[2][32+30].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+30].info_i__max_slave__  = 0.023000000;
slave_timing[2][32+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][32+30].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+30].t_rxd1[0][1] = 2334ns;
slave_timing[2][32+30].t_rxd1[1][0] = 2216ns;
slave_timing[2][32+30].t_rxd1[0][2] = 1781ns;
slave_timing[2][32+30].t_rxd1[2][0] = 2853ns;
slave_timing[2][32+30].t_rxd2[0][2] = 3590ns;
slave_timing[2][32+30].t_rxd2[2][0] = 2209ns;
slave_timing[2][32+30].t_rxd2[1][2] = 3250ns;
slave_timing[2][32+30].t_rxd2[2][1] = 2815ns;

slave_timing[2][32+31].info_corner          = 2;
slave_timing[2][32+31].info_temp__j__       = 125;
slave_timing[2][32+31].info_i__quite_rec__  = 0.040000000;
slave_timing[2][32+31].info_dtr__ib__       = 1;
slave_timing[2][32+31].info_i__offset_rec__ = 0.000000000;
slave_timing[2][32+31].info_i__max_slave__  = 0.025000000;
slave_timing[2][32+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][32+31].info_r__dsi_bus__    = 5.000;

slave_timing[2][32+31].t_rxd1[0][1] = 2256ns;
slave_timing[2][32+31].t_rxd1[1][0] = 2277ns;
slave_timing[2][32+31].t_rxd1[0][2] = 1733ns;
slave_timing[2][32+31].t_rxd1[2][0] = 2969ns;
slave_timing[2][32+31].t_rxd2[0][2] = 3312ns;
slave_timing[2][32+31].t_rxd2[2][0] = 2394ns;
slave_timing[2][32+31].t_rxd2[1][2] = 2906ns;
slave_timing[2][32+31].t_rxd2[2][1] = 3216ns;

/* ###   interface instances   ###################################################### */

ring_buffer_registers_BUF_VALID_COUNT_if ring_buffer_registers_BUF_VALID_COUNT (); 
ring_buffer_registers_BUF_FREE_if ring_buffer_registers_BUF_FREE (); 
ring_buffer_registers_BUF_READ_POINTER_if ring_buffer_registers_BUF_READ_POINTER (); 
ring_buffer_registers_BUF_WRITE_POINTER_if ring_buffer_registers_BUF_WRITE_POINTER (); 
ring_buffer_registers_BUF_VALID_POINTER_if ring_buffer_registers_BUF_VALID_POINTER (); 


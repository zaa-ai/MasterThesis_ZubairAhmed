
slave_timing[2][0].info_corner          = 1;
slave_timing[2][0].info_temp__j__       = 125;
slave_timing[2][0].info_i__quite_rec__  = 0.006000000;
slave_timing[2][0].info_dtr__ib__       = -1;
slave_timing[2][0].info_i__offset_rec__ = 0.000000000;
slave_timing[2][0].info_i__max_slave__  = 0.023000000;
slave_timing[2][0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][0].info_r__dsi_bus__    = 5.000;

slave_timing[2][0].t_rxd1[0][1] = 2196ns;
slave_timing[2][0].t_rxd1[1][0] = 2196ns;
slave_timing[2][0].t_rxd1[0][2] = 1662ns;
slave_timing[2][0].t_rxd1[2][0] = 2665ns;
slave_timing[2][0].t_rxd2[0][2] = 2617ns;
slave_timing[2][0].t_rxd2[2][0] = 1654ns;
slave_timing[2][0].t_rxd2[1][2] = 2172ns;
slave_timing[2][0].t_rxd2[2][1] = 2159ns;

slave_timing[2][1].info_corner          = 1;
slave_timing[2][1].info_temp__j__       = 125;
slave_timing[2][1].info_i__quite_rec__  = 0.006000000;
slave_timing[2][1].info_dtr__ib__       = -1;
slave_timing[2][1].info_i__offset_rec__ = 0.000000000;
slave_timing[2][1].info_i__max_slave__  = 0.025000000;
slave_timing[2][1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][1].info_r__dsi_bus__    = 5.000;

slave_timing[2][1].t_rxd1[0][1] = 2103ns;
slave_timing[2][1].t_rxd1[1][0] = 2265ns;
slave_timing[2][1].t_rxd1[0][2] = 1615ns;
slave_timing[2][1].t_rxd1[2][0] = 2707ns;
slave_timing[2][1].t_rxd2[0][2] = 2471ns;
slave_timing[2][1].t_rxd2[2][0] = 1762ns;
slave_timing[2][1].t_rxd2[1][2] = 1941ns;
slave_timing[2][1].t_rxd2[2][1] = 2390ns;

slave_timing[2][2].info_corner          = 1;
slave_timing[2][2].info_temp__j__       = 125;
slave_timing[2][2].info_i__quite_rec__  = 0.006000000;
slave_timing[2][2].info_dtr__ib__       = 1;
slave_timing[2][2].info_i__offset_rec__ = 0.000000000;
slave_timing[2][2].info_i__max_slave__  = 0.023000000;
slave_timing[2][2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][2].info_r__dsi_bus__    = 5.000;

slave_timing[2][2].t_rxd1[0][1] = 2269ns;
slave_timing[2][2].t_rxd1[1][0] = 2128ns;
slave_timing[2][2].t_rxd1[0][2] = 1699ns;
slave_timing[2][2].t_rxd1[2][0] = 2605ns;
slave_timing[2][2].t_rxd2[0][2] = 2765ns;
slave_timing[2][2].t_rxd2[2][0] = 1524ns;
slave_timing[2][2].t_rxd2[1][2] = 2396ns;
slave_timing[2][2].t_rxd2[2][1] = 1963ns;

slave_timing[2][3].info_corner          = 1;
slave_timing[2][3].info_temp__j__       = 125;
slave_timing[2][3].info_i__quite_rec__  = 0.006000000;
slave_timing[2][3].info_dtr__ib__       = 1;
slave_timing[2][3].info_i__offset_rec__ = 0.000000000;
slave_timing[2][3].info_i__max_slave__  = 0.025000000;
slave_timing[2][3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][3].info_r__dsi_bus__    = 5.000;

slave_timing[2][3].t_rxd1[0][1] = 2173ns;
slave_timing[2][3].t_rxd1[1][0] = 2200ns;
slave_timing[2][3].t_rxd1[0][2] = 1649ns;
slave_timing[2][3].t_rxd1[2][0] = 2650ns;
slave_timing[2][3].t_rxd2[0][2] = 2601ns;
slave_timing[2][3].t_rxd2[2][0] = 1667ns;
slave_timing[2][3].t_rxd2[1][2] = 2136ns;
slave_timing[2][3].t_rxd2[2][1] = 2189ns;

slave_timing[2][4].info_corner          = 1;
slave_timing[2][4].info_temp__j__       = 125;
slave_timing[2][4].info_i__quite_rec__  = 0.006000000;
slave_timing[2][4].info_dtr__ib__       = -1;
slave_timing[2][4].info_i__offset_rec__ = 0.000000000;
slave_timing[2][4].info_i__max_slave__  = 0.023000000;
slave_timing[2][4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][4].info_r__dsi_bus__    = 5.000;

slave_timing[2][4].t_rxd1[0][1] = 2381ns;
slave_timing[2][4].t_rxd1[1][0] = 2348ns;
slave_timing[2][4].t_rxd1[0][2] = 1825ns;
slave_timing[2][4].t_rxd1[2][0] = 2810ns;
slave_timing[2][4].t_rxd2[0][2] = 2654ns;
slave_timing[2][4].t_rxd2[2][0] = 1684ns;
slave_timing[2][4].t_rxd2[1][2] = 2199ns;
slave_timing[2][4].t_rxd2[2][1] = 2175ns;

slave_timing[2][5].info_corner          = 1;
slave_timing[2][5].info_temp__j__       = 125;
slave_timing[2][5].info_i__quite_rec__  = 0.006000000;
slave_timing[2][5].info_dtr__ib__       = -1;
slave_timing[2][5].info_i__offset_rec__ = 0.000000000;
slave_timing[2][5].info_i__max_slave__  = 0.025000000;
slave_timing[2][5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][5].info_r__dsi_bus__    = 5.000;

slave_timing[2][5].t_rxd1[0][1] = 2290ns;
slave_timing[2][5].t_rxd1[1][0] = 2423ns;
slave_timing[2][5].t_rxd1[0][2] = 1773ns;
slave_timing[2][5].t_rxd1[2][0] = 2849ns;
slave_timing[2][5].t_rxd2[0][2] = 2508ns;
slave_timing[2][5].t_rxd2[2][0] = 1799ns;
slave_timing[2][5].t_rxd2[1][2] = 1963ns;
slave_timing[2][5].t_rxd2[2][1] = 2426ns;

slave_timing[2][6].info_corner          = 1;
slave_timing[2][6].info_temp__j__       = 125;
slave_timing[2][6].info_i__quite_rec__  = 0.006000000;
slave_timing[2][6].info_dtr__ib__       = 1;
slave_timing[2][6].info_i__offset_rec__ = 0.000000000;
slave_timing[2][6].info_i__max_slave__  = 0.023000000;
slave_timing[2][6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][6].info_r__dsi_bus__    = 5.000;

slave_timing[2][6].t_rxd1[0][1] = 2469ns;
slave_timing[2][6].t_rxd1[1][0] = 2285ns;
slave_timing[2][6].t_rxd1[0][2] = 1863ns;
slave_timing[2][6].t_rxd1[2][0] = 2750ns;
slave_timing[2][6].t_rxd2[0][2] = 2803ns;
slave_timing[2][6].t_rxd2[2][0] = 1566ns;
slave_timing[2][6].t_rxd2[1][2] = 2419ns;
slave_timing[2][6].t_rxd2[2][1] = 2006ns;

slave_timing[2][7].info_corner          = 1;
slave_timing[2][7].info_temp__j__       = 125;
slave_timing[2][7].info_i__quite_rec__  = 0.006000000;
slave_timing[2][7].info_dtr__ib__       = 1;
slave_timing[2][7].info_i__offset_rec__ = 0.000000000;
slave_timing[2][7].info_i__max_slave__  = 0.025000000;
slave_timing[2][7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][7].info_r__dsi_bus__    = 5.000;

slave_timing[2][7].t_rxd1[0][1] = 2374ns;
slave_timing[2][7].t_rxd1[1][0] = 2348ns;
slave_timing[2][7].t_rxd1[0][2] = 1810ns;
slave_timing[2][7].t_rxd1[2][0] = 2793ns;
slave_timing[2][7].t_rxd2[0][2] = 2631ns;
slave_timing[2][7].t_rxd2[2][0] = 1697ns;
slave_timing[2][7].t_rxd2[1][2] = 2170ns;
slave_timing[2][7].t_rxd2[2][1] = 2228ns;

slave_timing[2][8].info_corner          = 1;
slave_timing[2][8].info_temp__j__       = 125;
slave_timing[2][8].info_i__quite_rec__  = 0.003000000;
slave_timing[2][8].info_dtr__ib__       = -1;
slave_timing[2][8].info_i__offset_rec__ = 0.000000000;
slave_timing[2][8].info_i__max_slave__  = 0.023000000;
slave_timing[2][8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][8].info_r__dsi_bus__    = 5.000;

slave_timing[2][8].t_rxd1[0][1] = 2155ns;
slave_timing[2][8].t_rxd1[1][0] = 2197ns;
slave_timing[2][8].t_rxd1[0][2] = 1643ns;
slave_timing[2][8].t_rxd1[2][0] = 2652ns;
slave_timing[2][8].t_rxd2[0][2] = 2598ns;
slave_timing[2][8].t_rxd2[2][0] = 1663ns;
slave_timing[2][8].t_rxd2[1][2] = 2133ns;
slave_timing[2][8].t_rxd2[2][1] = 2186ns;

slave_timing[2][9].info_corner          = 1;
slave_timing[2][9].info_temp__j__       = 125;
slave_timing[2][9].info_i__quite_rec__  = 0.003000000;
slave_timing[2][9].info_dtr__ib__       = -1;
slave_timing[2][9].info_i__offset_rec__ = 0.000000000;
slave_timing[2][9].info_i__max_slave__  = 0.025000000;
slave_timing[2][9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][9].info_r__dsi_bus__    = 5.000;

slave_timing[2][9].t_rxd1[0][1] = 2076ns;
slave_timing[2][9].t_rxd1[1][0] = 2261ns;
slave_timing[2][9].t_rxd1[0][2] = 1595ns;
slave_timing[2][9].t_rxd1[2][0] = 2698ns;
slave_timing[2][9].t_rxd2[0][2] = 2454ns;
slave_timing[2][9].t_rxd2[2][0] = 1771ns;
slave_timing[2][9].t_rxd2[1][2] = 1917ns;
slave_timing[2][9].t_rxd2[2][1] = 2413ns;

slave_timing[2][10].info_corner          = 1;
slave_timing[2][10].info_temp__j__       = 125;
slave_timing[2][10].info_i__quite_rec__  = 0.003000000;
slave_timing[2][10].info_dtr__ib__       = 1;
slave_timing[2][10].info_i__offset_rec__ = 0.000000000;
slave_timing[2][10].info_i__max_slave__  = 0.023000000;
slave_timing[2][10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][10].info_r__dsi_bus__    = 5.000;

slave_timing[2][10].t_rxd1[0][1] = 2227ns;
slave_timing[2][10].t_rxd1[1][0] = 2123ns;
slave_timing[2][10].t_rxd1[0][2] = 1670ns;
slave_timing[2][10].t_rxd1[2][0] = 2602ns;
slave_timing[2][10].t_rxd2[0][2] = 2742ns;
slave_timing[2][10].t_rxd2[2][0] = 1538ns;
slave_timing[2][10].t_rxd2[1][2] = 2367ns;
slave_timing[2][10].t_rxd2[2][1] = 1978ns;

slave_timing[2][11].info_corner          = 1;
slave_timing[2][11].info_temp__j__       = 125;
slave_timing[2][11].info_i__quite_rec__  = 0.003000000;
slave_timing[2][11].info_dtr__ib__       = 1;
slave_timing[2][11].info_i__offset_rec__ = 0.000000000;
slave_timing[2][11].info_i__max_slave__  = 0.025000000;
slave_timing[2][11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][11].info_r__dsi_bus__    = 5.000;

slave_timing[2][11].t_rxd1[0][1] = 2136ns;
slave_timing[2][11].t_rxd1[1][0] = 2178ns;
slave_timing[2][11].t_rxd1[0][2] = 1622ns;
slave_timing[2][11].t_rxd1[2][0] = 2641ns;
slave_timing[2][11].t_rxd2[0][2] = 2571ns;
slave_timing[2][11].t_rxd2[2][0] = 1666ns;
slave_timing[2][11].t_rxd2[1][2] = 2105ns;
slave_timing[2][11].t_rxd2[2][1] = 2210ns;

slave_timing[2][12].info_corner          = 1;
slave_timing[2][12].info_temp__j__       = 125;
slave_timing[2][12].info_i__quite_rec__  = 0.003000000;
slave_timing[2][12].info_dtr__ib__       = -1;
slave_timing[2][12].info_i__offset_rec__ = 0.000000000;
slave_timing[2][12].info_i__max_slave__  = 0.023000000;
slave_timing[2][12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][12].info_r__dsi_bus__    = 5.000;

slave_timing[2][12].t_rxd1[0][1] = 2362ns;
slave_timing[2][12].t_rxd1[1][0] = 2346ns;
slave_timing[2][12].t_rxd1[0][2] = 1813ns;
slave_timing[2][12].t_rxd1[2][0] = 2801ns;
slave_timing[2][12].t_rxd2[0][2] = 2633ns;
slave_timing[2][12].t_rxd2[2][0] = 1693ns;
slave_timing[2][12].t_rxd2[1][2] = 2171ns;
slave_timing[2][12].t_rxd2[2][1] = 2207ns;

slave_timing[2][13].info_corner          = 1;
slave_timing[2][13].info_temp__j__       = 125;
slave_timing[2][13].info_i__quite_rec__  = 0.003000000;
slave_timing[2][13].info_dtr__ib__       = -1;
slave_timing[2][13].info_i__offset_rec__ = 0.000000000;
slave_timing[2][13].info_i__max_slave__  = 0.025000000;
slave_timing[2][13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][13].info_r__dsi_bus__    = 5.000;

slave_timing[2][13].t_rxd1[0][1] = 2271ns;
slave_timing[2][13].t_rxd1[1][0] = 2411ns;
slave_timing[2][13].t_rxd1[0][2] = 1761ns;
slave_timing[2][13].t_rxd1[2][0] = 2840ns;
slave_timing[2][13].t_rxd2[0][2] = 2489ns;
slave_timing[2][13].t_rxd2[2][0] = 1798ns;
slave_timing[2][13].t_rxd2[1][2] = 1944ns;
slave_timing[2][13].t_rxd2[2][1] = 2433ns;

slave_timing[2][14].info_corner          = 1;
slave_timing[2][14].info_temp__j__       = 125;
slave_timing[2][14].info_i__quite_rec__  = 0.003000000;
slave_timing[2][14].info_dtr__ib__       = 1;
slave_timing[2][14].info_i__offset_rec__ = 0.000000000;
slave_timing[2][14].info_i__max_slave__  = 0.023000000;
slave_timing[2][14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][14].info_r__dsi_bus__    = 5.000;

slave_timing[2][14].t_rxd1[0][1] = 2423ns;
slave_timing[2][14].t_rxd1[1][0] = 2267ns;
slave_timing[2][14].t_rxd1[0][2] = 1843ns;
slave_timing[2][14].t_rxd1[2][0] = 2741ns;
slave_timing[2][14].t_rxd2[0][2] = 2770ns;
slave_timing[2][14].t_rxd2[2][0] = 1569ns;
slave_timing[2][14].t_rxd2[1][2] = 2380ns;
slave_timing[2][14].t_rxd2[2][1] = 2016ns;

slave_timing[2][15].info_corner          = 1;
slave_timing[2][15].info_temp__j__       = 125;
slave_timing[2][15].info_i__quite_rec__  = 0.003000000;
slave_timing[2][15].info_dtr__ib__       = 1;
slave_timing[2][15].info_i__offset_rec__ = 0.000000000;
slave_timing[2][15].info_i__max_slave__  = 0.025000000;
slave_timing[2][15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][15].info_r__dsi_bus__    = 5.000;

slave_timing[2][15].t_rxd1[0][1] = 2331ns;
slave_timing[2][15].t_rxd1[1][0] = 2343ns;
slave_timing[2][15].t_rxd1[0][2] = 1790ns;
slave_timing[2][15].t_rxd1[2][0] = 2783ns;
slave_timing[2][15].t_rxd2[0][2] = 2597ns;
slave_timing[2][15].t_rxd2[2][0] = 1698ns;
slave_timing[2][15].t_rxd2[1][2] = 2131ns;
slave_timing[2][15].t_rxd2[2][1] = 2232ns;

slave_timing[2][16].info_corner          = 1;
slave_timing[2][16].info_temp__j__       = 125;
slave_timing[2][16].info_i__quite_rec__  = 0.000000000;
slave_timing[2][16].info_dtr__ib__       = -1;
slave_timing[2][16].info_i__offset_rec__ = 0.000000000;
slave_timing[2][16].info_i__max_slave__  = 0.023000000;
slave_timing[2][16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][16].info_r__dsi_bus__    = 5.000;

slave_timing[2][16].t_rxd1[0][1] = 2146ns;
slave_timing[2][16].t_rxd1[1][0] = 2171ns;
slave_timing[2][16].t_rxd1[0][2] = 1611ns;
slave_timing[2][16].t_rxd1[2][0] = 2632ns;
slave_timing[2][16].t_rxd2[0][2] = 2571ns;
slave_timing[2][16].t_rxd2[2][0] = 1638ns;
slave_timing[2][16].t_rxd2[1][2] = 2141ns;
slave_timing[2][16].t_rxd2[2][1] = 2164ns;

slave_timing[2][17].info_corner          = 1;
slave_timing[2][17].info_temp__j__       = 125;
slave_timing[2][17].info_i__quite_rec__  = 0.000000000;
slave_timing[2][17].info_dtr__ib__       = -1;
slave_timing[2][17].info_i__offset_rec__ = 0.000000000;
slave_timing[2][17].info_i__max_slave__  = 0.025000000;
slave_timing[2][17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][17].info_r__dsi_bus__    = 5.000;

slave_timing[2][17].t_rxd1[0][1] = 2065ns;
slave_timing[2][17].t_rxd1[1][0] = 2244ns;
slave_timing[2][17].t_rxd1[0][2] = 1577ns;
slave_timing[2][17].t_rxd1[2][0] = 2667ns;
slave_timing[2][17].t_rxd2[0][2] = 2443ns;
slave_timing[2][17].t_rxd2[2][0] = 1752ns;
slave_timing[2][17].t_rxd2[1][2] = 1930ns;
slave_timing[2][17].t_rxd2[2][1] = 2382ns;

slave_timing[2][18].info_corner          = 1;
slave_timing[2][18].info_temp__j__       = 125;
slave_timing[2][18].info_i__quite_rec__  = 0.000000000;
slave_timing[2][18].info_dtr__ib__       = 1;
slave_timing[2][18].info_i__offset_rec__ = 0.000000000;
slave_timing[2][18].info_i__max_slave__  = 0.023000000;
slave_timing[2][18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][18].info_r__dsi_bus__    = 5.000;

slave_timing[2][18].t_rxd1[0][1] = 2234ns;
slave_timing[2][18].t_rxd1[1][0] = 2055ns;
slave_timing[2][18].t_rxd1[0][2] = 1672ns;
slave_timing[2][18].t_rxd1[2][0] = 2550ns;
slave_timing[2][18].t_rxd2[0][2] = 2764ns;
slave_timing[2][18].t_rxd2[2][0] = 1489ns;
slave_timing[2][18].t_rxd2[1][2] = 2392ns;
slave_timing[2][18].t_rxd2[2][1] = 1907ns;

slave_timing[2][19].info_corner          = 1;
slave_timing[2][19].info_temp__j__       = 125;
slave_timing[2][19].info_i__quite_rec__  = 0.000000000;
slave_timing[2][19].info_dtr__ib__       = 1;
slave_timing[2][19].info_i__offset_rec__ = 0.000000000;
slave_timing[2][19].info_i__max_slave__  = 0.025000000;
slave_timing[2][19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][19].info_r__dsi_bus__    = 5.000;

slave_timing[2][19].t_rxd1[0][1] = 2152ns;
slave_timing[2][19].t_rxd1[1][0] = 2135ns;
slave_timing[2][19].t_rxd1[0][2] = 1622ns;
slave_timing[2][19].t_rxd1[2][0] = 2592ns;
slave_timing[2][19].t_rxd2[0][2] = 2574ns;
slave_timing[2][19].t_rxd2[2][0] = 1628ns;
slave_timing[2][19].t_rxd2[1][2] = 2136ns;
slave_timing[2][19].t_rxd2[2][1] = 2135ns;

slave_timing[2][20].info_corner          = 1;
slave_timing[2][20].info_temp__j__       = 125;
slave_timing[2][20].info_i__quite_rec__  = 0.000000000;
slave_timing[2][20].info_dtr__ib__       = -1;
slave_timing[2][20].info_i__offset_rec__ = 0.000000000;
slave_timing[2][20].info_i__max_slave__  = 0.023000000;
slave_timing[2][20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][20].info_r__dsi_bus__    = 5.000;

slave_timing[2][20].t_rxd1[0][1] = 2370ns;
slave_timing[2][20].t_rxd1[1][0] = 2316ns;
slave_timing[2][20].t_rxd1[0][2] = 1814ns;
slave_timing[2][20].t_rxd1[2][0] = 2771ns;
slave_timing[2][20].t_rxd2[0][2] = 2626ns;
slave_timing[2][20].t_rxd2[2][0] = 1669ns;
slave_timing[2][20].t_rxd2[1][2] = 2175ns;
slave_timing[2][20].t_rxd2[2][1] = 2179ns;

slave_timing[2][21].info_corner          = 1;
slave_timing[2][21].info_temp__j__       = 125;
slave_timing[2][21].info_i__quite_rec__  = 0.000000000;
slave_timing[2][21].info_dtr__ib__       = -1;
slave_timing[2][21].info_i__offset_rec__ = 0.000000000;
slave_timing[2][21].info_i__max_slave__  = 0.025000000;
slave_timing[2][21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][21].info_r__dsi_bus__    = 5.000;

slave_timing[2][21].t_rxd1[0][1] = 2276ns;
slave_timing[2][21].t_rxd1[1][0] = 2384ns;
slave_timing[2][21].t_rxd1[0][2] = 1764ns;
slave_timing[2][21].t_rxd1[2][0] = 2810ns;
slave_timing[2][21].t_rxd2[0][2] = 2481ns;
slave_timing[2][21].t_rxd2[2][0] = 1782ns;
slave_timing[2][21].t_rxd2[1][2] = 1941ns;
slave_timing[2][21].t_rxd2[2][1] = 2406ns;

slave_timing[2][22].info_corner          = 1;
slave_timing[2][22].info_temp__j__       = 125;
slave_timing[2][22].info_i__quite_rec__  = 0.000000000;
slave_timing[2][22].info_dtr__ib__       = 1;
slave_timing[2][22].info_i__offset_rec__ = 0.000000000;
slave_timing[2][22].info_i__max_slave__  = 0.023000000;
slave_timing[2][22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][22].info_r__dsi_bus__    = 5.000;

slave_timing[2][22].t_rxd1[0][1] = 2458ns;
slave_timing[2][22].t_rxd1[1][0] = 2233ns;
slave_timing[2][22].t_rxd1[0][2] = 1859ns;
slave_timing[2][22].t_rxd1[2][0] = 2693ns;
slave_timing[2][22].t_rxd2[0][2] = 2790ns;
slave_timing[2][22].t_rxd2[2][0] = 1516ns;
slave_timing[2][22].t_rxd2[1][2] = 2431ns;
slave_timing[2][22].t_rxd2[2][1] = 1913ns;

slave_timing[2][23].info_corner          = 1;
slave_timing[2][23].info_temp__j__       = 125;
slave_timing[2][23].info_i__quite_rec__  = 0.000000000;
slave_timing[2][23].info_dtr__ib__       = 1;
slave_timing[2][23].info_i__offset_rec__ = 0.000000000;
slave_timing[2][23].info_i__max_slave__  = 0.025000000;
slave_timing[2][23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][23].info_r__dsi_bus__    = 5.000;

slave_timing[2][23].t_rxd1[0][1] = 2363ns;
slave_timing[2][23].t_rxd1[1][0] = 2296ns;
slave_timing[2][23].t_rxd1[0][2] = 1806ns;
slave_timing[2][23].t_rxd1[2][0] = 2733ns;
slave_timing[2][23].t_rxd2[0][2] = 2605ns;
slave_timing[2][23].t_rxd2[2][0] = 1649ns;
slave_timing[2][23].t_rxd2[1][2] = 2169ns;
slave_timing[2][23].t_rxd2[2][1] = 2156ns;

slave_timing[2][24].info_corner          = 1;
slave_timing[2][24].info_temp__j__       = 125;
slave_timing[2][24].info_i__quite_rec__  = 0.040000000;
slave_timing[2][24].info_dtr__ib__       = -1;
slave_timing[2][24].info_i__offset_rec__ = 0.000000000;
slave_timing[2][24].info_i__max_slave__  = 0.023000000;
slave_timing[2][24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][24].info_r__dsi_bus__    = 5.000;

slave_timing[2][24].t_rxd1[0][1] = 2173ns;
slave_timing[2][24].t_rxd1[1][0] = 2244ns;
slave_timing[2][24].t_rxd1[0][2] = 1642ns;
slave_timing[2][24].t_rxd1[2][0] = 2681ns;
slave_timing[2][24].t_rxd2[0][2] = 2611ns;
slave_timing[2][24].t_rxd2[2][0] = 1675ns;
slave_timing[2][24].t_rxd2[1][2] = 2178ns;
slave_timing[2][24].t_rxd2[2][1] = 2188ns;

slave_timing[2][25].info_corner          = 1;
slave_timing[2][25].info_temp__j__       = 125;
slave_timing[2][25].info_i__quite_rec__  = 0.040000000;
slave_timing[2][25].info_dtr__ib__       = -1;
slave_timing[2][25].info_i__offset_rec__ = 0.000000000;
slave_timing[2][25].info_i__max_slave__  = 0.025000000;
slave_timing[2][25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][25].info_r__dsi_bus__    = 5.000;

slave_timing[2][25].t_rxd1[0][1] = 2091ns;
slave_timing[2][25].t_rxd1[1][0] = 2299ns;
slave_timing[2][25].t_rxd1[0][2] = 1596ns;
slave_timing[2][25].t_rxd1[2][0] = 2724ns;
slave_timing[2][25].t_rxd2[0][2] = 2462ns;
slave_timing[2][25].t_rxd2[2][0] = 1776ns;
slave_timing[2][25].t_rxd2[1][2] = 1919ns;
slave_timing[2][25].t_rxd2[2][1] = 2439ns;

slave_timing[2][26].info_corner          = 1;
slave_timing[2][26].info_temp__j__       = 125;
slave_timing[2][26].info_i__quite_rec__  = 0.040000000;
slave_timing[2][26].info_dtr__ib__       = 1;
slave_timing[2][26].info_i__offset_rec__ = 0.000000000;
slave_timing[2][26].info_i__max_slave__  = 0.023000000;
slave_timing[2][26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][26].info_r__dsi_bus__    = 5.000;

slave_timing[2][26].t_rxd1[0][1] = 2249ns;
slave_timing[2][26].t_rxd1[1][0] = 2133ns;
slave_timing[2][26].t_rxd1[0][2] = 1690ns;
slave_timing[2][26].t_rxd1[2][0] = 2621ns;
slave_timing[2][26].t_rxd2[0][2] = 2762ns;
slave_timing[2][26].t_rxd2[2][0] = 1554ns;
slave_timing[2][26].t_rxd2[1][2] = 2366ns;
slave_timing[2][26].t_rxd2[2][1] = 2002ns;

slave_timing[2][27].info_corner          = 1;
slave_timing[2][27].info_temp__j__       = 125;
slave_timing[2][27].info_i__quite_rec__  = 0.040000000;
slave_timing[2][27].info_dtr__ib__       = 1;
slave_timing[2][27].info_i__offset_rec__ = 0.000000000;
slave_timing[2][27].info_i__max_slave__  = 0.025000000;
slave_timing[2][27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[2][27].info_r__dsi_bus__    = 5.000;

slave_timing[2][27].t_rxd1[0][1] = 2162ns;
slave_timing[2][27].t_rxd1[1][0] = 2211ns;
slave_timing[2][27].t_rxd1[0][2] = 1628ns;
slave_timing[2][27].t_rxd1[2][0] = 2665ns;
slave_timing[2][27].t_rxd2[0][2] = 2585ns;
slave_timing[2][27].t_rxd2[2][0] = 1683ns;
slave_timing[2][27].t_rxd2[1][2] = 2113ns;
slave_timing[2][27].t_rxd2[2][1] = 2199ns;

slave_timing[2][28].info_corner          = 1;
slave_timing[2][28].info_temp__j__       = 125;
slave_timing[2][28].info_i__quite_rec__  = 0.040000000;
slave_timing[2][28].info_dtr__ib__       = -1;
slave_timing[2][28].info_i__offset_rec__ = 0.000000000;
slave_timing[2][28].info_i__max_slave__  = 0.023000000;
slave_timing[2][28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][28].info_r__dsi_bus__    = 5.000;

slave_timing[2][28].t_rxd1[0][1] = 2259ns;
slave_timing[2][28].t_rxd1[1][0] = 2336ns;
slave_timing[2][28].t_rxd1[0][2] = 1741ns;
slave_timing[2][28].t_rxd1[2][0] = 2764ns;
slave_timing[2][28].t_rxd2[0][2] = 2642ns;
slave_timing[2][28].t_rxd2[2][0] = 1712ns;
slave_timing[2][28].t_rxd2[1][2] = 2220ns;
slave_timing[2][28].t_rxd2[2][1] = 2207ns;

slave_timing[2][29].info_corner          = 1;
slave_timing[2][29].info_temp__j__       = 125;
slave_timing[2][29].info_i__quite_rec__  = 0.040000000;
slave_timing[2][29].info_dtr__ib__       = -1;
slave_timing[2][29].info_i__offset_rec__ = 0.000000000;
slave_timing[2][29].info_i__max_slave__  = 0.025000000;
slave_timing[2][29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][29].info_r__dsi_bus__    = 5.000;

slave_timing[2][29].t_rxd1[0][1] = 2187ns;
slave_timing[2][29].t_rxd1[1][0] = 2395ns;
slave_timing[2][29].t_rxd1[0][2] = 1693ns;
slave_timing[2][29].t_rxd1[2][0] = 2816ns;
slave_timing[2][29].t_rxd2[0][2] = 2504ns;
slave_timing[2][29].t_rxd2[2][0] = 1811ns;
slave_timing[2][29].t_rxd2[1][2] = 1977ns;
slave_timing[2][29].t_rxd2[2][1] = 2435ns;

slave_timing[2][30].info_corner          = 1;
slave_timing[2][30].info_temp__j__       = 125;
slave_timing[2][30].info_i__quite_rec__  = 0.040000000;
slave_timing[2][30].info_dtr__ib__       = 1;
slave_timing[2][30].info_i__offset_rec__ = 0.000000000;
slave_timing[2][30].info_i__max_slave__  = 0.023000000;
slave_timing[2][30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][30].info_r__dsi_bus__    = 5.000;

slave_timing[2][30].t_rxd1[0][1] = 2353ns;
slave_timing[2][30].t_rxd1[1][0] = 2233ns;
slave_timing[2][30].t_rxd1[0][2] = 1785ns;
slave_timing[2][30].t_rxd1[2][0] = 2713ns;
slave_timing[2][30].t_rxd2[0][2] = 2792ns;
slave_timing[2][30].t_rxd2[2][0] = 1590ns;
slave_timing[2][30].t_rxd2[1][2] = 2399ns;
slave_timing[2][30].t_rxd2[2][1] = 2037ns;

slave_timing[2][31].info_corner          = 1;
slave_timing[2][31].info_temp__j__       = 125;
slave_timing[2][31].info_i__quite_rec__  = 0.040000000;
slave_timing[2][31].info_dtr__ib__       = 1;
slave_timing[2][31].info_i__offset_rec__ = 0.000000000;
slave_timing[2][31].info_i__max_slave__  = 0.025000000;
slave_timing[2][31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[2][31].info_r__dsi_bus__    = 5.000;

slave_timing[2][31].t_rxd1[0][1] = 2262ns;
slave_timing[2][31].t_rxd1[1][0] = 2307ns;
slave_timing[2][31].t_rxd1[0][2] = 1732ns;
slave_timing[2][31].t_rxd1[2][0] = 2755ns;
slave_timing[2][31].t_rxd2[0][2] = 2628ns;
slave_timing[2][31].t_rxd2[2][0] = 1702ns;
slave_timing[2][31].t_rxd2[1][2] = 2151ns;
slave_timing[2][31].t_rxd2[2][1] = 2257ns;

/* ###   interface instances   ###################################################### */

JTAG_standard_registers_JTAG_ID_if JTAG_standard_registers_JTAG_ID (); 
JTAG_standard_registers_JTAG_BYPASS_if JTAG_standard_registers_JTAG_BYPASS (); 



slave_timing[3][224+0].info_corner          = 4;
slave_timing[3][224+0].info_temp__j__       = -40;
slave_timing[3][224+0].info_i__quite_rec__  = 0.006000000;
slave_timing[3][224+0].info_dtr__ib__       = -1;
slave_timing[3][224+0].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+0].info_i__max_slave__  = 0.023000000;
slave_timing[3][224+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][224+0].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+0].t_rxd1[0][1] = 2796ns;
slave_timing[3][224+0].t_rxd1[1][0] = 2749ns;
slave_timing[3][224+0].t_rxd1[0][2] = 2088ns;
slave_timing[3][224+0].t_rxd1[2][0] = 3363ns;
slave_timing[3][224+0].t_rxd2[0][2] = 3378ns;
slave_timing[3][224+0].t_rxd2[2][0] = 2054ns;
slave_timing[3][224+0].t_rxd2[1][2] = 2790ns;
slave_timing[3][224+0].t_rxd2[2][1] = 2730ns;

slave_timing[3][224+1].info_corner          = 4;
slave_timing[3][224+1].info_temp__j__       = -40;
slave_timing[3][224+1].info_i__quite_rec__  = 0.006000000;
slave_timing[3][224+1].info_dtr__ib__       = -1;
slave_timing[3][224+1].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+1].info_i__max_slave__  = 0.025000000;
slave_timing[3][224+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][224+1].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+1].t_rxd1[0][1] = 2687ns;
slave_timing[3][224+1].t_rxd1[1][0] = 2835ns;
slave_timing[3][224+1].t_rxd1[0][2] = 2024ns;
slave_timing[3][224+1].t_rxd1[2][0] = 3420ns;
slave_timing[3][224+1].t_rxd2[0][2] = 3182ns;
slave_timing[3][224+1].t_rxd2[2][0] = 2206ns;
slave_timing[3][224+1].t_rxd2[1][2] = 2527ns;
slave_timing[3][224+1].t_rxd2[2][1] = 2976ns;

slave_timing[3][224+2].info_corner          = 4;
slave_timing[3][224+2].info_temp__j__       = -40;
slave_timing[3][224+2].info_i__quite_rec__  = 0.006000000;
slave_timing[3][224+2].info_dtr__ib__       = 1;
slave_timing[3][224+2].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+2].info_i__max_slave__  = 0.023000000;
slave_timing[3][224+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][224+2].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+2].t_rxd1[0][1] = 2862ns;
slave_timing[3][224+2].t_rxd1[1][0] = 2699ns;
slave_timing[3][224+2].t_rxd1[0][2] = 2120ns;
slave_timing[3][224+2].t_rxd1[2][0] = 3331ns;
slave_timing[3][224+2].t_rxd2[0][2] = 3529ns;
slave_timing[3][224+2].t_rxd2[2][0] = 1943ns;
slave_timing[3][224+2].t_rxd2[1][2] = 3007ns;
slave_timing[3][224+2].t_rxd2[2][1] = 2538ns;

slave_timing[3][224+3].info_corner          = 4;
slave_timing[3][224+3].info_temp__j__       = -40;
slave_timing[3][224+3].info_i__quite_rec__  = 0.006000000;
slave_timing[3][224+3].info_dtr__ib__       = 1;
slave_timing[3][224+3].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+3].info_i__max_slave__  = 0.025000000;
slave_timing[3][224+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][224+3].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+3].t_rxd1[0][1] = 2747ns;
slave_timing[3][224+3].t_rxd1[1][0] = 2789ns;
slave_timing[3][224+3].t_rxd1[0][2] = 2057ns;
slave_timing[3][224+3].t_rxd1[2][0] = 3388ns;
slave_timing[3][224+3].t_rxd2[0][2] = 3301ns;
slave_timing[3][224+3].t_rxd2[2][0] = 2116ns;
slave_timing[3][224+3].t_rxd2[1][2] = 2668ns;
slave_timing[3][224+3].t_rxd2[2][1] = 2795ns;

slave_timing[3][224+4].info_corner          = 4;
slave_timing[3][224+4].info_temp__j__       = -40;
slave_timing[3][224+4].info_i__quite_rec__  = 0.006000000;
slave_timing[3][224+4].info_dtr__ib__       = -1;
slave_timing[3][224+4].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+4].info_i__max_slave__  = 0.023000000;
slave_timing[3][224+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][224+4].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+4].t_rxd1[0][1] = 2874ns;
slave_timing[3][224+4].t_rxd1[1][0] = 2821ns;
slave_timing[3][224+4].t_rxd1[0][2] = 2153ns;
slave_timing[3][224+4].t_rxd1[2][0] = 3432ns;
slave_timing[3][224+4].t_rxd2[0][2] = 3390ns;
slave_timing[3][224+4].t_rxd2[2][0] = 2068ns;
slave_timing[3][224+4].t_rxd2[1][2] = 2805ns;
slave_timing[3][224+4].t_rxd2[2][1] = 2734ns;

slave_timing[3][224+5].info_corner          = 4;
slave_timing[3][224+5].info_temp__j__       = -40;
slave_timing[3][224+5].info_i__quite_rec__  = 0.006000000;
slave_timing[3][224+5].info_dtr__ib__       = -1;
slave_timing[3][224+5].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+5].info_i__max_slave__  = 0.025000000;
slave_timing[3][224+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][224+5].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+5].t_rxd1[0][1] = 2762ns;
slave_timing[3][224+5].t_rxd1[1][0] = 2905ns;
slave_timing[3][224+5].t_rxd1[0][2] = 2086ns;
slave_timing[3][224+5].t_rxd1[2][0] = 3488ns;
slave_timing[3][224+5].t_rxd2[0][2] = 3197ns;
slave_timing[3][224+5].t_rxd2[2][0] = 2217ns;
slave_timing[3][224+5].t_rxd2[1][2] = 2505ns;
slave_timing[3][224+5].t_rxd2[2][1] = 3030ns;

slave_timing[3][224+6].info_corner          = 4;
slave_timing[3][224+6].info_temp__j__       = -40;
slave_timing[3][224+6].info_i__quite_rec__  = 0.006000000;
slave_timing[3][224+6].info_dtr__ib__       = 1;
slave_timing[3][224+6].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+6].info_i__max_slave__  = 0.023000000;
slave_timing[3][224+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][224+6].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+6].t_rxd1[0][1] = 2931ns;
slave_timing[3][224+6].t_rxd1[1][0] = 2768ns;
slave_timing[3][224+6].t_rxd1[0][2] = 2184ns;
slave_timing[3][224+6].t_rxd1[2][0] = 3396ns;
slave_timing[3][224+6].t_rxd2[0][2] = 3540ns;
slave_timing[3][224+6].t_rxd2[2][0] = 1954ns;
slave_timing[3][224+6].t_rxd2[1][2] = 3014ns;
slave_timing[3][224+6].t_rxd2[2][1] = 2516ns;

slave_timing[3][224+7].info_corner          = 4;
slave_timing[3][224+7].info_temp__j__       = -40;
slave_timing[3][224+7].info_i__quite_rec__  = 0.006000000;
slave_timing[3][224+7].info_dtr__ib__       = 1;
slave_timing[3][224+7].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+7].info_i__max_slave__  = 0.025000000;
slave_timing[3][224+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][224+7].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+7].t_rxd1[0][1] = 2812ns;
slave_timing[3][224+7].t_rxd1[1][0] = 2853ns;
slave_timing[3][224+7].t_rxd1[0][2] = 2119ns;
slave_timing[3][224+7].t_rxd1[2][0] = 3453ns;
slave_timing[3][224+7].t_rxd2[0][2] = 3313ns;
slave_timing[3][224+7].t_rxd2[2][0] = 2126ns;
slave_timing[3][224+7].t_rxd2[1][2] = 2684ns;
slave_timing[3][224+7].t_rxd2[2][1] = 2836ns;

slave_timing[3][224+8].info_corner          = 4;
slave_timing[3][224+8].info_temp__j__       = -40;
slave_timing[3][224+8].info_i__quite_rec__  = 0.003000000;
slave_timing[3][224+8].info_dtr__ib__       = -1;
slave_timing[3][224+8].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+8].info_i__max_slave__  = 0.023000000;
slave_timing[3][224+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][224+8].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+8].t_rxd1[0][1] = 2774ns;
slave_timing[3][224+8].t_rxd1[1][0] = 2767ns;
slave_timing[3][224+8].t_rxd1[0][2] = 2077ns;
slave_timing[3][224+8].t_rxd1[2][0] = 3377ns;
slave_timing[3][224+8].t_rxd2[0][2] = 3364ns;
slave_timing[3][224+8].t_rxd2[2][0] = 2062ns;
slave_timing[3][224+8].t_rxd2[1][2] = 2767ns;
slave_timing[3][224+8].t_rxd2[2][1] = 2705ns;

slave_timing[3][224+9].info_corner          = 4;
slave_timing[3][224+9].info_temp__j__       = -40;
slave_timing[3][224+9].info_i__quite_rec__  = 0.003000000;
slave_timing[3][224+9].info_dtr__ib__       = -1;
slave_timing[3][224+9].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+9].info_i__max_slave__  = 0.025000000;
slave_timing[3][224+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][224+9].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+9].t_rxd1[0][1] = 2671ns;
slave_timing[3][224+9].t_rxd1[1][0] = 2852ns;
slave_timing[3][224+9].t_rxd1[0][2] = 2011ns;
slave_timing[3][224+9].t_rxd1[2][0] = 3435ns;
slave_timing[3][224+9].t_rxd2[0][2] = 3169ns;
slave_timing[3][224+9].t_rxd2[2][0] = 2212ns;
slave_timing[3][224+9].t_rxd2[1][2] = 2475ns;
slave_timing[3][224+9].t_rxd2[2][1] = 3032ns;

slave_timing[3][224+10].info_corner          = 4;
slave_timing[3][224+10].info_temp__j__       = -40;
slave_timing[3][224+10].info_i__quite_rec__  = 0.003000000;
slave_timing[3][224+10].info_dtr__ib__       = 1;
slave_timing[3][224+10].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+10].info_i__max_slave__  = 0.023000000;
slave_timing[3][224+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][224+10].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+10].t_rxd1[0][1] = 2849ns;
slave_timing[3][224+10].t_rxd1[1][0] = 2708ns;
slave_timing[3][224+10].t_rxd1[0][2] = 2114ns;
slave_timing[3][224+10].t_rxd1[2][0] = 3339ns;
slave_timing[3][224+10].t_rxd2[0][2] = 3516ns;
slave_timing[3][224+10].t_rxd2[2][0] = 1948ns;
slave_timing[3][224+10].t_rxd2[1][2] = 2986ns;
slave_timing[3][224+10].t_rxd2[2][1] = 2557ns;

slave_timing[3][224+11].info_corner          = 4;
slave_timing[3][224+11].info_temp__j__       = -40;
slave_timing[3][224+11].info_i__quite_rec__  = 0.003000000;
slave_timing[3][224+11].info_dtr__ib__       = 1;
slave_timing[3][224+11].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+11].info_i__max_slave__  = 0.025000000;
slave_timing[3][224+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][224+11].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+11].t_rxd1[0][1] = 2735ns;
slave_timing[3][224+11].t_rxd1[1][0] = 2799ns;
slave_timing[3][224+11].t_rxd1[0][2] = 2049ns;
slave_timing[3][224+11].t_rxd1[2][0] = 3395ns;
slave_timing[3][224+11].t_rxd2[0][2] = 3290ns;
slave_timing[3][224+11].t_rxd2[2][0] = 2118ns;
slave_timing[3][224+11].t_rxd2[1][2] = 2656ns;
slave_timing[3][224+11].t_rxd2[2][1] = 2846ns;

slave_timing[3][224+12].info_corner          = 4;
slave_timing[3][224+12].info_temp__j__       = -40;
slave_timing[3][224+12].info_i__quite_rec__  = 0.003000000;
slave_timing[3][224+12].info_dtr__ib__       = -1;
slave_timing[3][224+12].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+12].info_i__max_slave__  = 0.023000000;
slave_timing[3][224+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][224+12].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+12].t_rxd1[0][1] = 2857ns;
slave_timing[3][224+12].t_rxd1[1][0] = 2839ns;
slave_timing[3][224+12].t_rxd1[0][2] = 2145ns;
slave_timing[3][224+12].t_rxd1[2][0] = 3448ns;
slave_timing[3][224+12].t_rxd2[0][2] = 3376ns;
slave_timing[3][224+12].t_rxd2[2][0] = 2076ns;
slave_timing[3][224+12].t_rxd2[1][2] = 2820ns;
slave_timing[3][224+12].t_rxd2[2][1] = 2715ns;

slave_timing[3][224+13].info_corner          = 4;
slave_timing[3][224+13].info_temp__j__       = -40;
slave_timing[3][224+13].info_i__quite_rec__  = 0.003000000;
slave_timing[3][224+13].info_dtr__ib__       = -1;
slave_timing[3][224+13].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+13].info_i__max_slave__  = 0.025000000;
slave_timing[3][224+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][224+13].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+13].t_rxd1[0][1] = 2746ns;
slave_timing[3][224+13].t_rxd1[1][0] = 2922ns;
slave_timing[3][224+13].t_rxd1[0][2] = 2085ns;
slave_timing[3][224+13].t_rxd1[2][0] = 3502ns;
slave_timing[3][224+13].t_rxd2[0][2] = 3185ns;
slave_timing[3][224+13].t_rxd2[2][0] = 2227ns;
slave_timing[3][224+13].t_rxd2[1][2] = 2482ns;
slave_timing[3][224+13].t_rxd2[2][1] = 3044ns;

slave_timing[3][224+14].info_corner          = 4;
slave_timing[3][224+14].info_temp__j__       = -40;
slave_timing[3][224+14].info_i__quite_rec__  = 0.003000000;
slave_timing[3][224+14].info_dtr__ib__       = 1;
slave_timing[3][224+14].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+14].info_i__max_slave__  = 0.023000000;
slave_timing[3][224+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][224+14].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+14].t_rxd1[0][1] = 2918ns;
slave_timing[3][224+14].t_rxd1[1][0] = 2779ns;
slave_timing[3][224+14].t_rxd1[0][2] = 2179ns;
slave_timing[3][224+14].t_rxd1[2][0] = 3401ns;
slave_timing[3][224+14].t_rxd2[0][2] = 3528ns;
slave_timing[3][224+14].t_rxd2[2][0] = 1954ns;
slave_timing[3][224+14].t_rxd2[1][2] = 2996ns;
slave_timing[3][224+14].t_rxd2[2][1] = 2560ns;

slave_timing[3][224+15].info_corner          = 4;
slave_timing[3][224+15].info_temp__j__       = -40;
slave_timing[3][224+15].info_i__quite_rec__  = 0.003000000;
slave_timing[3][224+15].info_dtr__ib__       = 1;
slave_timing[3][224+15].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+15].info_i__max_slave__  = 0.025000000;
slave_timing[3][224+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][224+15].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+15].t_rxd1[0][1] = 2804ns;
slave_timing[3][224+15].t_rxd1[1][0] = 2866ns;
slave_timing[3][224+15].t_rxd1[0][2] = 2110ns;
slave_timing[3][224+15].t_rxd1[2][0] = 3461ns;
slave_timing[3][224+15].t_rxd2[0][2] = 3300ns;
slave_timing[3][224+15].t_rxd2[2][0] = 2130ns;
slave_timing[3][224+15].t_rxd2[1][2] = 2670ns;
slave_timing[3][224+15].t_rxd2[2][1] = 2853ns;

slave_timing[3][224+16].info_corner          = 4;
slave_timing[3][224+16].info_temp__j__       = -40;
slave_timing[3][224+16].info_i__quite_rec__  = 0.000000000;
slave_timing[3][224+16].info_dtr__ib__       = -1;
slave_timing[3][224+16].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+16].info_i__max_slave__  = 0.023000000;
slave_timing[3][224+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][224+16].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+16].t_rxd1[0][1] = 2800ns;
slave_timing[3][224+16].t_rxd1[1][0] = 2750ns;
slave_timing[3][224+16].t_rxd1[0][2] = 2069ns;
slave_timing[3][224+16].t_rxd1[2][0] = 3363ns;
slave_timing[3][224+16].t_rxd2[0][2] = 3350ns;
slave_timing[3][224+16].t_rxd2[2][0] = 2052ns;
slave_timing[3][224+16].t_rxd2[1][2] = 2792ns;
slave_timing[3][224+16].t_rxd2[2][1] = 2731ns;

slave_timing[3][224+17].info_corner          = 4;
slave_timing[3][224+17].info_temp__j__       = -40;
slave_timing[3][224+17].info_i__quite_rec__  = 0.000000000;
slave_timing[3][224+17].info_dtr__ib__       = -1;
slave_timing[3][224+17].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+17].info_i__max_slave__  = 0.025000000;
slave_timing[3][224+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][224+17].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+17].t_rxd1[0][1] = 2692ns;
slave_timing[3][224+17].t_rxd1[1][0] = 2836ns;
slave_timing[3][224+17].t_rxd1[0][2] = 2004ns;
slave_timing[3][224+17].t_rxd1[2][0] = 3421ns;
slave_timing[3][224+17].t_rxd2[0][2] = 3161ns;
slave_timing[3][224+17].t_rxd2[2][0] = 2225ns;
slave_timing[3][224+17].t_rxd2[1][2] = 2492ns;
slave_timing[3][224+17].t_rxd2[2][1] = 3017ns;

slave_timing[3][224+18].info_corner          = 4;
slave_timing[3][224+18].info_temp__j__       = -40;
slave_timing[3][224+18].info_i__quite_rec__  = 0.000000000;
slave_timing[3][224+18].info_dtr__ib__       = 1;
slave_timing[3][224+18].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+18].info_i__max_slave__  = 0.023000000;
slave_timing[3][224+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][224+18].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+18].t_rxd1[0][1] = 2835ns;
slave_timing[3][224+18].t_rxd1[1][0] = 2733ns;
slave_timing[3][224+18].t_rxd1[0][2] = 2110ns;
slave_timing[3][224+18].t_rxd1[2][0] = 3354ns;
slave_timing[3][224+18].t_rxd2[0][2] = 3506ns;
slave_timing[3][224+18].t_rxd2[2][0] = 1959ns;
slave_timing[3][224+18].t_rxd2[1][2] = 2974ns;
slave_timing[3][224+18].t_rxd2[2][1] = 2565ns;

slave_timing[3][224+19].info_corner          = 4;
slave_timing[3][224+19].info_temp__j__       = -40;
slave_timing[3][224+19].info_i__quite_rec__  = 0.000000000;
slave_timing[3][224+19].info_dtr__ib__       = 1;
slave_timing[3][224+19].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+19].info_i__max_slave__  = 0.025000000;
slave_timing[3][224+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][224+19].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+19].t_rxd1[0][1] = 2720ns;
slave_timing[3][224+19].t_rxd1[1][0] = 2817ns;
slave_timing[3][224+19].t_rxd1[0][2] = 2044ns;
slave_timing[3][224+19].t_rxd1[2][0] = 3408ns;
slave_timing[3][224+19].t_rxd2[0][2] = 3281ns;
slave_timing[3][224+19].t_rxd2[2][0] = 2126ns;
slave_timing[3][224+19].t_rxd2[1][2] = 2643ns;
slave_timing[3][224+19].t_rxd2[2][1] = 2855ns;

slave_timing[3][224+20].info_corner          = 4;
slave_timing[3][224+20].info_temp__j__       = -40;
slave_timing[3][224+20].info_i__quite_rec__  = 0.000000000;
slave_timing[3][224+20].info_dtr__ib__       = -1;
slave_timing[3][224+20].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+20].info_i__max_slave__  = 0.023000000;
slave_timing[3][224+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][224+20].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+20].t_rxd1[0][1] = 2880ns;
slave_timing[3][224+20].t_rxd1[1][0] = 2818ns;
slave_timing[3][224+20].t_rxd1[0][2] = 2139ns;
slave_timing[3][224+20].t_rxd1[2][0] = 3430ns;
slave_timing[3][224+20].t_rxd2[0][2] = 3364ns;
slave_timing[3][224+20].t_rxd2[2][0] = 2067ns;
slave_timing[3][224+20].t_rxd2[1][2] = 2793ns;
slave_timing[3][224+20].t_rxd2[2][1] = 2735ns;

slave_timing[3][224+21].info_corner          = 4;
slave_timing[3][224+21].info_temp__j__       = -40;
slave_timing[3][224+21].info_i__quite_rec__  = 0.000000000;
slave_timing[3][224+21].info_dtr__ib__       = -1;
slave_timing[3][224+21].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+21].info_i__max_slave__  = 0.025000000;
slave_timing[3][224+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][224+21].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+21].t_rxd1[0][1] = 2768ns;
slave_timing[3][224+21].t_rxd1[1][0] = 2902ns;
slave_timing[3][224+21].t_rxd1[0][2] = 2075ns;
slave_timing[3][224+21].t_rxd1[2][0] = 3513ns;
slave_timing[3][224+21].t_rxd2[0][2] = 3172ns;
slave_timing[3][224+21].t_rxd2[2][0] = 2237ns;
slave_timing[3][224+21].t_rxd2[1][2] = 2504ns;
slave_timing[3][224+21].t_rxd2[2][1] = 3025ns;

slave_timing[3][224+22].info_corner          = 4;
slave_timing[3][224+22].info_temp__j__       = -40;
slave_timing[3][224+22].info_i__quite_rec__  = 0.000000000;
slave_timing[3][224+22].info_dtr__ib__       = 1;
slave_timing[3][224+22].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+22].info_i__max_slave__  = 0.023000000;
slave_timing[3][224+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][224+22].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+22].t_rxd1[0][1] = 2953ns;
slave_timing[3][224+22].t_rxd1[1][0] = 2752ns;
slave_timing[3][224+22].t_rxd1[0][2] = 2166ns;
slave_timing[3][224+22].t_rxd1[2][0] = 3414ns;
slave_timing[3][224+22].t_rxd2[0][2] = 3514ns;
slave_timing[3][224+22].t_rxd2[2][0] = 1965ns;
slave_timing[3][224+22].t_rxd2[1][2] = 3024ns;
slave_timing[3][224+22].t_rxd2[2][1] = 2534ns;

slave_timing[3][224+23].info_corner          = 4;
slave_timing[3][224+23].info_temp__j__       = -40;
slave_timing[3][224+23].info_i__quite_rec__  = 0.000000000;
slave_timing[3][224+23].info_dtr__ib__       = 1;
slave_timing[3][224+23].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+23].info_i__max_slave__  = 0.025000000;
slave_timing[3][224+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][224+23].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+23].t_rxd1[0][1] = 2791ns;
slave_timing[3][224+23].t_rxd1[1][0] = 2879ns;
slave_timing[3][224+23].t_rxd1[0][2] = 2110ns;
slave_timing[3][224+23].t_rxd1[2][0] = 3468ns;
slave_timing[3][224+23].t_rxd2[0][2] = 3294ns;
slave_timing[3][224+23].t_rxd2[2][0] = 2136ns;
slave_timing[3][224+23].t_rxd2[1][2] = 2657ns;
slave_timing[3][224+23].t_rxd2[2][1] = 2864ns;

slave_timing[3][224+24].info_corner          = 4;
slave_timing[3][224+24].info_temp__j__       = -40;
slave_timing[3][224+24].info_i__quite_rec__  = 0.040000000;
slave_timing[3][224+24].info_dtr__ib__       = -1;
slave_timing[3][224+24].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+24].info_i__max_slave__  = 0.023000000;
slave_timing[3][224+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][224+24].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+24].t_rxd1[0][1] = 2796ns;
slave_timing[3][224+24].t_rxd1[1][0] = 2731ns;
slave_timing[3][224+24].t_rxd1[0][2] = 2061ns;
slave_timing[3][224+24].t_rxd1[2][0] = 3375ns;
slave_timing[3][224+24].t_rxd2[0][2] = 3360ns;
slave_timing[3][224+24].t_rxd2[2][0] = 2071ns;
slave_timing[3][224+24].t_rxd2[1][2] = 2799ns;
slave_timing[3][224+24].t_rxd2[2][1] = 2718ns;

slave_timing[3][224+25].info_corner          = 4;
slave_timing[3][224+25].info_temp__j__       = -40;
slave_timing[3][224+25].info_i__quite_rec__  = 0.040000000;
slave_timing[3][224+25].info_dtr__ib__       = -1;
slave_timing[3][224+25].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+25].info_i__max_slave__  = 0.025000000;
slave_timing[3][224+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][224+25].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+25].t_rxd1[0][1] = 2650ns;
slave_timing[3][224+25].t_rxd1[1][0] = 2853ns;
slave_timing[3][224+25].t_rxd1[0][2] = 1999ns;
slave_timing[3][224+25].t_rxd1[2][0] = 3429ns;
slave_timing[3][224+25].t_rxd2[0][2] = 3167ns;
slave_timing[3][224+25].t_rxd2[2][0] = 2219ns;
slave_timing[3][224+25].t_rxd2[1][2] = 2504ns;
slave_timing[3][224+25].t_rxd2[2][1] = 3005ns;

slave_timing[3][224+26].info_corner          = 4;
slave_timing[3][224+26].info_temp__j__       = -40;
slave_timing[3][224+26].info_i__quite_rec__  = 0.040000000;
slave_timing[3][224+26].info_dtr__ib__       = 1;
slave_timing[3][224+26].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+26].info_i__max_slave__  = 0.023000000;
slave_timing[3][224+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][224+26].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+26].t_rxd1[0][1] = 2845ns;
slave_timing[3][224+26].t_rxd1[1][0] = 2697ns;
slave_timing[3][224+26].t_rxd1[0][2] = 2110ns;
slave_timing[3][224+26].t_rxd1[2][0] = 3330ns;
slave_timing[3][224+26].t_rxd2[0][2] = 3524ns;
slave_timing[3][224+26].t_rxd2[2][0] = 1945ns;
slave_timing[3][224+26].t_rxd2[1][2] = 2998ns;
slave_timing[3][224+26].t_rxd2[2][1] = 2549ns;

slave_timing[3][224+27].info_corner          = 4;
slave_timing[3][224+27].info_temp__j__       = -40;
slave_timing[3][224+27].info_i__quite_rec__  = 0.040000000;
slave_timing[3][224+27].info_dtr__ib__       = 1;
slave_timing[3][224+27].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+27].info_i__max_slave__  = 0.025000000;
slave_timing[3][224+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][224+27].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+27].t_rxd1[0][1] = 2734ns;
slave_timing[3][224+27].t_rxd1[1][0] = 2787ns;
slave_timing[3][224+27].t_rxd1[0][2] = 2044ns;
slave_timing[3][224+27].t_rxd1[2][0] = 3385ns;
slave_timing[3][224+27].t_rxd2[0][2] = 3296ns;
slave_timing[3][224+27].t_rxd2[2][0] = 2117ns;
slave_timing[3][224+27].t_rxd2[1][2] = 2668ns;
slave_timing[3][224+27].t_rxd2[2][1] = 2842ns;

slave_timing[3][224+28].info_corner          = 4;
slave_timing[3][224+28].info_temp__j__       = -40;
slave_timing[3][224+28].info_i__quite_rec__  = 0.040000000;
slave_timing[3][224+28].info_dtr__ib__       = -1;
slave_timing[3][224+28].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+28].info_i__max_slave__  = 0.023000000;
slave_timing[3][224+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][224+28].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+28].t_rxd1[0][1] = 2832ns;
slave_timing[3][224+28].t_rxd1[1][0] = 2766ns;
slave_timing[3][224+28].t_rxd1[0][2] = 2091ns;
slave_timing[3][224+28].t_rxd1[2][0] = 3410ns;
slave_timing[3][224+28].t_rxd2[0][2] = 3372ns;
slave_timing[3][224+28].t_rxd2[2][0] = 2084ns;
slave_timing[3][224+28].t_rxd2[1][2] = 2818ns;
slave_timing[3][224+28].t_rxd2[2][1] = 2731ns;

slave_timing[3][224+29].info_corner          = 4;
slave_timing[3][224+29].info_temp__j__       = -40;
slave_timing[3][224+29].info_i__quite_rec__  = 0.040000000;
slave_timing[3][224+29].info_dtr__ib__       = -1;
slave_timing[3][224+29].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+29].info_i__max_slave__  = 0.025000000;
slave_timing[3][224+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][224+29].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+29].t_rxd1[0][1] = 2684ns;
slave_timing[3][224+29].t_rxd1[1][0] = 2891ns;
slave_timing[3][224+29].t_rxd1[0][2] = 2031ns;
slave_timing[3][224+29].t_rxd1[2][0] = 3463ns;
slave_timing[3][224+29].t_rxd2[0][2] = 3183ns;
slave_timing[3][224+29].t_rxd2[2][0] = 2238ns;
slave_timing[3][224+29].t_rxd2[1][2] = 2483ns;
slave_timing[3][224+29].t_rxd2[2][1] = 3056ns;

slave_timing[3][224+30].info_corner          = 4;
slave_timing[3][224+30].info_temp__j__       = -40;
slave_timing[3][224+30].info_i__quite_rec__  = 0.040000000;
slave_timing[3][224+30].info_dtr__ib__       = 1;
slave_timing[3][224+30].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+30].info_i__max_slave__  = 0.023000000;
slave_timing[3][224+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][224+30].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+30].t_rxd1[0][1] = 2879ns;
slave_timing[3][224+30].t_rxd1[1][0] = 2733ns;
slave_timing[3][224+30].t_rxd1[0][2] = 2142ns;
slave_timing[3][224+30].t_rxd1[2][0] = 3360ns;
slave_timing[3][224+30].t_rxd2[0][2] = 3537ns;
slave_timing[3][224+30].t_rxd2[2][0] = 1956ns;
slave_timing[3][224+30].t_rxd2[1][2] = 3014ns;
slave_timing[3][224+30].t_rxd2[2][1] = 2562ns;

slave_timing[3][224+31].info_corner          = 4;
slave_timing[3][224+31].info_temp__j__       = -40;
slave_timing[3][224+31].info_i__quite_rec__  = 0.040000000;
slave_timing[3][224+31].info_dtr__ib__       = 1;
slave_timing[3][224+31].info_i__offset_rec__ = 0.000000000;
slave_timing[3][224+31].info_i__max_slave__  = 0.025000000;
slave_timing[3][224+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][224+31].info_r__dsi_bus__    = 5.000;

slave_timing[3][224+31].t_rxd1[0][1] = 2762ns;
slave_timing[3][224+31].t_rxd1[1][0] = 2818ns;
slave_timing[3][224+31].t_rxd1[0][2] = 2077ns;
slave_timing[3][224+31].t_rxd1[2][0] = 3416ns;
slave_timing[3][224+31].t_rxd2[0][2] = 3311ns;
slave_timing[3][224+31].t_rxd2[2][0] = 2128ns;
slave_timing[3][224+31].t_rxd2[1][2] = 2679ns;
slave_timing[3][224+31].t_rxd2[2][1] = 2853ns;

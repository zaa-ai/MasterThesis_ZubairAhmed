
slave_timing[0][0].info_corner          = 0;
slave_timing[0][0].info_temp__j__       = 25;
slave_timing[0][0].info_i__quite_rec__  = 0.006000000;
slave_timing[0][0].info_dtr__ib__       = -1;
slave_timing[0][0].info_i__offset_rec__ = -0.001000000;
slave_timing[0][0].info_i__max_slave__  = 0.021000000;
slave_timing[0][0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][0].info_r__dsi_bus__    = 5.000;

slave_timing[0][0].t_rxd1[0][1] = 1514ns;
slave_timing[0][0].t_rxd1[1][0] = 1044ns;
slave_timing[0][0].t_rxd1[0][2] = 983ns;
slave_timing[0][0].t_rxd1[2][0] = 1356ns;
slave_timing[0][0].t_rxd2[0][2] = 1783ns;
slave_timing[0][0].t_rxd2[2][0] = 813ns;
slave_timing[0][0].t_rxd2[1][2] = 1535ns;
slave_timing[0][0].t_rxd2[2][1] = 1047ns;

slave_timing[0][1].info_corner          = 0;
slave_timing[0][1].info_temp__j__       = 25;
slave_timing[0][1].info_i__quite_rec__  = 0.006000000;
slave_timing[0][1].info_dtr__ib__       = -1;
slave_timing[0][1].info_i__offset_rec__ = 0.001000000;
slave_timing[0][1].info_i__max_slave__  = 0.021000000;
slave_timing[0][1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][1].info_r__dsi_bus__    = 5.000;

slave_timing[0][1].t_rxd1[0][1] = 1224ns;
slave_timing[0][1].t_rxd1[1][0] = 1249ns;
slave_timing[0][1].t_rxd1[0][2] = 891ns;
slave_timing[0][1].t_rxd1[2][0] = 1531ns;
slave_timing[0][1].t_rxd2[0][2] = 1507ns;
slave_timing[0][1].t_rxd2[2][0] = 910ns;
slave_timing[0][1].t_rxd2[1][2] = 1234ns;
slave_timing[0][1].t_rxd2[2][1] = 1251ns;

slave_timing[0][2].info_corner          = 0;
slave_timing[0][2].info_temp__j__       = 25;
slave_timing[0][2].info_i__quite_rec__  = 0.006000000;
slave_timing[0][2].info_dtr__ib__       = -1;
slave_timing[0][2].info_i__offset_rec__ = -0.001000000;
slave_timing[0][2].info_i__max_slave__  = 0.027000000;
slave_timing[0][2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][2].info_r__dsi_bus__    = 5.000;

slave_timing[0][2].t_rxd1[0][1] = 1233ns;
slave_timing[0][2].t_rxd1[1][0] = 1162ns;
slave_timing[0][2].t_rxd1[0][2] = 893ns;
slave_timing[0][2].t_rxd1[2][0] = 1453ns;
slave_timing[0][2].t_rxd2[0][2] = 1318ns;
slave_timing[0][2].t_rxd2[2][0] = 978ns;
slave_timing[0][2].t_rxd2[1][2] = 1005ns;
slave_timing[0][2].t_rxd2[2][1] = 1484ns;

slave_timing[0][3].info_corner          = 0;
slave_timing[0][3].info_temp__j__       = 25;
slave_timing[0][3].info_i__quite_rec__  = 0.006000000;
slave_timing[0][3].info_dtr__ib__       = -1;
slave_timing[0][3].info_i__offset_rec__ = 0.001000000;
slave_timing[0][3].info_i__max_slave__  = 0.027000000;
slave_timing[0][3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][3].info_r__dsi_bus__    = 5.000;

slave_timing[0][3].t_rxd1[0][1] = 1086ns;
slave_timing[0][3].t_rxd1[1][0] = 1328ns;
slave_timing[0][3].t_rxd1[0][2] = 816ns;
slave_timing[0][3].t_rxd1[2][0] = 1602ns;
slave_timing[0][3].t_rxd2[0][2] = 1220ns;
slave_timing[0][3].t_rxd2[2][0] = 1042ns;
slave_timing[0][3].t_rxd2[1][2] = 872ns;
slave_timing[0][3].t_rxd2[2][1] = 1910ns;

slave_timing[0][4].info_corner          = 0;
slave_timing[0][4].info_temp__j__       = 25;
slave_timing[0][4].info_i__quite_rec__  = 0.006000000;
slave_timing[0][4].info_dtr__ib__       = 1;
slave_timing[0][4].info_i__offset_rec__ = -0.001000000;
slave_timing[0][4].info_i__max_slave__  = 0.021000000;
slave_timing[0][4].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][4].info_r__dsi_bus__    = 5.000;

slave_timing[0][4].t_rxd1[0][1] = 1620ns;
slave_timing[0][4].t_rxd1[1][0] = 1017ns;
slave_timing[0][4].t_rxd1[0][2] = 1005ns;
slave_timing[0][4].t_rxd1[2][0] = 1334ns;
slave_timing[0][4].t_rxd2[0][2] = 2122ns;
slave_timing[0][4].t_rxd2[2][0] = 762ns;
slave_timing[0][4].t_rxd2[1][2] = 1882ns;
slave_timing[0][4].t_rxd2[2][1] = 955ns;

slave_timing[0][5].info_corner          = 0;
slave_timing[0][5].info_temp__j__       = 25;
slave_timing[0][5].info_i__quite_rec__  = 0.006000000;
slave_timing[0][5].info_dtr__ib__       = 1;
slave_timing[0][5].info_i__offset_rec__ = 0.001000000;
slave_timing[0][5].info_i__max_slave__  = 0.021000000;
slave_timing[0][5].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][5].info_r__dsi_bus__    = 5.000;

slave_timing[0][5].t_rxd1[0][1] = 1278ns;
slave_timing[0][5].t_rxd1[1][0] = 1214ns;
slave_timing[0][5].t_rxd1[0][2] = 912ns;
slave_timing[0][5].t_rxd1[2][0] = 1500ns;
slave_timing[0][5].t_rxd2[0][2] = 1644ns;
slave_timing[0][5].t_rxd2[2][0] = 864ns;
slave_timing[0][5].t_rxd2[1][2] = 1386ns;
slave_timing[0][5].t_rxd2[2][1] = 1144ns;

slave_timing[0][6].info_corner          = 0;
slave_timing[0][6].info_temp__j__       = 25;
slave_timing[0][6].info_i__quite_rec__  = 0.006000000;
slave_timing[0][6].info_dtr__ib__       = 1;
slave_timing[0][6].info_i__offset_rec__ = -0.001000000;
slave_timing[0][6].info_i__max_slave__  = 0.027000000;
slave_timing[0][6].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][6].info_r__dsi_bus__    = 5.000;

slave_timing[0][6].t_rxd1[0][1] = 1273ns;
slave_timing[0][6].t_rxd1[1][0] = 1138ns;
slave_timing[0][6].t_rxd1[0][2] = 909ns;
slave_timing[0][6].t_rxd1[2][0] = 1431ns;
slave_timing[0][6].t_rxd2[0][2] = 1383ns;
slave_timing[0][6].t_rxd2[2][0] = 943ns;
slave_timing[0][6].t_rxd2[1][2] = 1091ns;
slave_timing[0][6].t_rxd2[2][1] = 1354ns;

slave_timing[0][7].info_corner          = 0;
slave_timing[0][7].info_temp__j__       = 25;
slave_timing[0][7].info_i__quite_rec__  = 0.006000000;
slave_timing[0][7].info_dtr__ib__       = 1;
slave_timing[0][7].info_i__offset_rec__ = 0.001000000;
slave_timing[0][7].info_i__max_slave__  = 0.027000000;
slave_timing[0][7].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][7].info_r__dsi_bus__    = 5.000;

slave_timing[0][7].t_rxd1[0][1] = 1122ns;
slave_timing[0][7].t_rxd1[1][0] = 1296ns;
slave_timing[0][7].t_rxd1[0][2] = 834ns;
slave_timing[0][7].t_rxd1[2][0] = 1593ns;
slave_timing[0][7].t_rxd2[0][2] = 1273ns;
slave_timing[0][7].t_rxd2[2][0] = 1015ns;
slave_timing[0][7].t_rxd2[1][2] = 960ns;
slave_timing[0][7].t_rxd2[2][1] = 1626ns;

slave_timing[0][8].info_corner          = 0;
slave_timing[0][8].info_temp__j__       = 25;
slave_timing[0][8].info_i__quite_rec__  = 0.006000000;
slave_timing[0][8].info_dtr__ib__       = -1;
slave_timing[0][8].info_i__offset_rec__ = -0.001000000;
slave_timing[0][8].info_i__max_slave__  = 0.021000000;
slave_timing[0][8].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][8].info_r__dsi_bus__    = 5.000;

slave_timing[0][8].t_rxd1[0][1] = 1801ns;
slave_timing[0][8].t_rxd1[1][0] = 1246ns;
slave_timing[0][8].t_rxd1[0][2] = 1177ns;
slave_timing[0][8].t_rxd1[2][0] = 1619ns;
slave_timing[0][8].t_rxd2[0][2] = 2113ns;
slave_timing[0][8].t_rxd2[2][0] = 971ns;
slave_timing[0][8].t_rxd2[1][2] = 1824ns;
slave_timing[0][8].t_rxd2[2][1] = 1246ns;

slave_timing[0][9].info_corner          = 0;
slave_timing[0][9].info_temp__j__       = 25;
slave_timing[0][9].info_i__quite_rec__  = 0.006000000;
slave_timing[0][9].info_dtr__ib__       = -1;
slave_timing[0][9].info_i__offset_rec__ = 0.001000000;
slave_timing[0][9].info_i__max_slave__  = 0.021000000;
slave_timing[0][9].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][9].info_r__dsi_bus__    = 5.000;

slave_timing[0][9].t_rxd1[0][1] = 1458ns;
slave_timing[0][9].t_rxd1[1][0] = 1492ns;
slave_timing[0][9].t_rxd1[0][2] = 1064ns;
slave_timing[0][9].t_rxd1[2][0] = 1823ns;
slave_timing[0][9].t_rxd2[0][2] = 1797ns;
slave_timing[0][9].t_rxd2[2][0] = 1085ns;
slave_timing[0][9].t_rxd2[1][2] = 1472ns;
slave_timing[0][9].t_rxd2[2][1] = 1495ns;

slave_timing[0][10].info_corner          = 0;
slave_timing[0][10].info_temp__j__       = 25;
slave_timing[0][10].info_i__quite_rec__  = 0.006000000;
slave_timing[0][10].info_dtr__ib__       = -1;
slave_timing[0][10].info_i__offset_rec__ = -0.001000000;
slave_timing[0][10].info_i__max_slave__  = 0.027000000;
slave_timing[0][10].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][10].info_r__dsi_bus__    = 5.000;

slave_timing[0][10].t_rxd1[0][1] = 1470ns;
slave_timing[0][10].t_rxd1[1][0] = 1390ns;
slave_timing[0][10].t_rxd1[0][2] = 1065ns;
slave_timing[0][10].t_rxd1[2][0] = 1734ns;
slave_timing[0][10].t_rxd2[0][2] = 1574ns;
slave_timing[0][10].t_rxd2[2][0] = 1168ns;
slave_timing[0][10].t_rxd2[1][2] = 1198ns;
slave_timing[0][10].t_rxd2[2][1] = 1769ns;

slave_timing[0][11].info_corner          = 0;
slave_timing[0][11].info_temp__j__       = 25;
slave_timing[0][11].info_i__quite_rec__  = 0.006000000;
slave_timing[0][11].info_dtr__ib__       = -1;
slave_timing[0][11].info_i__offset_rec__ = 0.001000000;
slave_timing[0][11].info_i__max_slave__  = 0.027000000;
slave_timing[0][11].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][11].info_r__dsi_bus__    = 5.000;

slave_timing[0][11].t_rxd1[0][1] = 1275ns;
slave_timing[0][11].t_rxd1[1][0] = 1614ns;
slave_timing[0][11].t_rxd1[0][2] = 977ns;
slave_timing[0][11].t_rxd1[2][0] = 1932ns;
slave_timing[0][11].t_rxd2[0][2] = 1459ns;
slave_timing[0][11].t_rxd2[2][0] = 1254ns;
slave_timing[0][11].t_rxd2[1][2] = 1026ns;
slave_timing[0][11].t_rxd2[2][1] = 2346ns;

slave_timing[0][12].info_corner          = 0;
slave_timing[0][12].info_temp__j__       = 25;
slave_timing[0][12].info_i__quite_rec__  = 0.006000000;
slave_timing[0][12].info_dtr__ib__       = 1;
slave_timing[0][12].info_i__offset_rec__ = -0.001000000;
slave_timing[0][12].info_i__max_slave__  = 0.021000000;
slave_timing[0][12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][12].info_r__dsi_bus__    = 5.000;

slave_timing[0][12].t_rxd1[0][1] = 1921ns;
slave_timing[0][12].t_rxd1[1][0] = 1211ns;
slave_timing[0][12].t_rxd1[0][2] = 1198ns;
slave_timing[0][12].t_rxd1[2][0] = 1594ns;
slave_timing[0][12].t_rxd2[0][2] = 2484ns;
slave_timing[0][12].t_rxd2[2][0] = 910ns;
slave_timing[0][12].t_rxd2[1][2] = 2219ns;
slave_timing[0][12].t_rxd2[2][1] = 1139ns;

slave_timing[0][13].info_corner          = 0;
slave_timing[0][13].info_temp__j__       = 25;
slave_timing[0][13].info_i__quite_rec__  = 0.006000000;
slave_timing[0][13].info_dtr__ib__       = 1;
slave_timing[0][13].info_i__offset_rec__ = 0.001000000;
slave_timing[0][13].info_i__max_slave__  = 0.021000000;
slave_timing[0][13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][13].info_r__dsi_bus__    = 5.000;

slave_timing[0][13].t_rxd1[0][1] = 1523ns;
slave_timing[0][13].t_rxd1[1][0] = 1447ns;
slave_timing[0][13].t_rxd1[0][2] = 1091ns;
slave_timing[0][13].t_rxd1[2][0] = 1788ns;
slave_timing[0][13].t_rxd2[0][2] = 1954ns;
slave_timing[0][13].t_rxd2[2][0] = 1032ns;
slave_timing[0][13].t_rxd2[1][2] = 1651ns;
slave_timing[0][13].t_rxd2[2][1] = 1363ns;

slave_timing[0][14].info_corner          = 0;
slave_timing[0][14].info_temp__j__       = 25;
slave_timing[0][14].info_i__quite_rec__  = 0.006000000;
slave_timing[0][14].info_dtr__ib__       = 1;
slave_timing[0][14].info_i__offset_rec__ = -0.001000000;
slave_timing[0][14].info_i__max_slave__  = 0.027000000;
slave_timing[0][14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][14].info_r__dsi_bus__    = 5.000;

slave_timing[0][14].t_rxd1[0][1] = 1520ns;
slave_timing[0][14].t_rxd1[1][0] = 1359ns;
slave_timing[0][14].t_rxd1[0][2] = 1084ns;
slave_timing[0][14].t_rxd1[2][0] = 1711ns;
slave_timing[0][14].t_rxd2[0][2] = 1652ns;
slave_timing[0][14].t_rxd2[2][0] = 1127ns;
slave_timing[0][14].t_rxd2[1][2] = 1301ns;
slave_timing[0][14].t_rxd2[2][1] = 1618ns;

slave_timing[0][15].info_corner          = 0;
slave_timing[0][15].info_temp__j__       = 25;
slave_timing[0][15].info_i__quite_rec__  = 0.006000000;
slave_timing[0][15].info_dtr__ib__       = 1;
slave_timing[0][15].info_i__offset_rec__ = 0.001000000;
slave_timing[0][15].info_i__max_slave__  = 0.027000000;
slave_timing[0][15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][15].info_r__dsi_bus__    = 5.000;

slave_timing[0][15].t_rxd1[0][1] = 1339ns;
slave_timing[0][15].t_rxd1[1][0] = 1551ns;
slave_timing[0][15].t_rxd1[0][2] = 999ns;
slave_timing[0][15].t_rxd1[2][0] = 1874ns;
slave_timing[0][15].t_rxd2[0][2] = 1523ns;
slave_timing[0][15].t_rxd2[2][0] = 1202ns;
slave_timing[0][15].t_rxd2[1][2] = 1143ns;
slave_timing[0][15].t_rxd2[2][1] = 1931ns;

slave_timing[0][16].info_corner          = 0;
slave_timing[0][16].info_temp__j__       = 25;
slave_timing[0][16].info_i__quite_rec__  = 0.003000000;
slave_timing[0][16].info_dtr__ib__       = -1;
slave_timing[0][16].info_i__offset_rec__ = -0.001000000;
slave_timing[0][16].info_i__max_slave__  = 0.021000000;
slave_timing[0][16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][16].info_r__dsi_bus__    = 5.000;

slave_timing[0][16].t_rxd1[0][1] = 1498ns;
slave_timing[0][16].t_rxd1[1][0] = 1047ns;
slave_timing[0][16].t_rxd1[0][2] = 980ns;
slave_timing[0][16].t_rxd1[2][0] = 1359ns;
slave_timing[0][16].t_rxd2[0][2] = 1768ns;
slave_timing[0][16].t_rxd2[2][0] = 817ns;
slave_timing[0][16].t_rxd2[1][2] = 1517ns;
slave_timing[0][16].t_rxd2[2][1] = 1054ns;

slave_timing[0][17].info_corner          = 0;
slave_timing[0][17].info_temp__j__       = 25;
slave_timing[0][17].info_i__quite_rec__  = 0.003000000;
slave_timing[0][17].info_dtr__ib__       = -1;
slave_timing[0][17].info_i__offset_rec__ = 0.001000000;
slave_timing[0][17].info_i__max_slave__  = 0.021000000;
slave_timing[0][17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][17].info_r__dsi_bus__    = 5.000;

slave_timing[0][17].t_rxd1[0][1] = 1213ns;
slave_timing[0][17].t_rxd1[1][0] = 1253ns;
slave_timing[0][17].t_rxd1[0][2] = 887ns;
slave_timing[0][17].t_rxd1[2][0] = 1533ns;
slave_timing[0][17].t_rxd2[0][2] = 1497ns;
slave_timing[0][17].t_rxd2[2][0] = 911ns;
slave_timing[0][17].t_rxd2[1][2] = 1228ns;
slave_timing[0][17].t_rxd2[2][1] = 1260ns;

slave_timing[0][18].info_corner          = 0;
slave_timing[0][18].info_temp__j__       = 25;
slave_timing[0][18].info_i__quite_rec__  = 0.003000000;
slave_timing[0][18].info_dtr__ib__       = -1;
slave_timing[0][18].info_i__offset_rec__ = -0.001000000;
slave_timing[0][18].info_i__max_slave__  = 0.027000000;
slave_timing[0][18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][18].info_r__dsi_bus__    = 5.000;

slave_timing[0][18].t_rxd1[0][1] = 1225ns;
slave_timing[0][18].t_rxd1[1][0] = 1163ns;
slave_timing[0][18].t_rxd1[0][2] = 898ns;
slave_timing[0][18].t_rxd1[2][0] = 1442ns;
slave_timing[0][18].t_rxd2[0][2] = 1323ns;
slave_timing[0][18].t_rxd2[2][0] = 974ns;
slave_timing[0][18].t_rxd2[1][2] = 998ns;
slave_timing[0][18].t_rxd2[2][1] = 1494ns;

slave_timing[0][19].info_corner          = 0;
slave_timing[0][19].info_temp__j__       = 25;
slave_timing[0][19].info_i__quite_rec__  = 0.003000000;
slave_timing[0][19].info_dtr__ib__       = -1;
slave_timing[0][19].info_i__offset_rec__ = 0.001000000;
slave_timing[0][19].info_i__max_slave__  = 0.027000000;
slave_timing[0][19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][19].info_r__dsi_bus__    = 5.000;

slave_timing[0][19].t_rxd1[0][1] = 1064ns;
slave_timing[0][19].t_rxd1[1][0] = 1356ns;
slave_timing[0][19].t_rxd1[0][2] = 815ns;
slave_timing[0][19].t_rxd1[2][0] = 1626ns;
slave_timing[0][19].t_rxd2[0][2] = 1216ns;
slave_timing[0][19].t_rxd2[2][0] = 1051ns;
slave_timing[0][19].t_rxd2[1][2] = 850ns;
slave_timing[0][19].t_rxd2[2][1] = 2034ns;

slave_timing[0][20].info_corner          = 0;
slave_timing[0][20].info_temp__j__       = 25;
slave_timing[0][20].info_i__quite_rec__  = 0.003000000;
slave_timing[0][20].info_dtr__ib__       = 1;
slave_timing[0][20].info_i__offset_rec__ = -0.001000000;
slave_timing[0][20].info_i__max_slave__  = 0.021000000;
slave_timing[0][20].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][20].info_r__dsi_bus__    = 5.000;

slave_timing[0][20].t_rxd1[0][1] = 1598ns;
slave_timing[0][20].t_rxd1[1][0] = 1020ns;
slave_timing[0][20].t_rxd1[0][2] = 1002ns;
slave_timing[0][20].t_rxd1[2][0] = 1337ns;
slave_timing[0][20].t_rxd2[0][2] = 2089ns;
slave_timing[0][20].t_rxd2[2][0] = 766ns;
slave_timing[0][20].t_rxd2[1][2] = 1847ns;
slave_timing[0][20].t_rxd2[2][1] = 963ns;

slave_timing[0][21].info_corner          = 0;
slave_timing[0][21].info_temp__j__       = 25;
slave_timing[0][21].info_i__quite_rec__  = 0.003000000;
slave_timing[0][21].info_dtr__ib__       = 1;
slave_timing[0][21].info_i__offset_rec__ = 0.001000000;
slave_timing[0][21].info_i__max_slave__  = 0.021000000;
slave_timing[0][21].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][21].info_r__dsi_bus__    = 5.000;

slave_timing[0][21].t_rxd1[0][1] = 1268ns;
slave_timing[0][21].t_rxd1[1][0] = 1218ns;
slave_timing[0][21].t_rxd1[0][2] = 910ns;
slave_timing[0][21].t_rxd1[2][0] = 1504ns;
slave_timing[0][21].t_rxd2[0][2] = 1632ns;
slave_timing[0][21].t_rxd2[2][0] = 867ns;
slave_timing[0][21].t_rxd2[1][2] = 1374ns;
slave_timing[0][21].t_rxd2[2][1] = 1153ns;

slave_timing[0][22].info_corner          = 0;
slave_timing[0][22].info_temp__j__       = 25;
slave_timing[0][22].info_i__quite_rec__  = 0.003000000;
slave_timing[0][22].info_dtr__ib__       = 1;
slave_timing[0][22].info_i__offset_rec__ = -0.001000000;
slave_timing[0][22].info_i__max_slave__  = 0.027000000;
slave_timing[0][22].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][22].info_r__dsi_bus__    = 5.000;

slave_timing[0][22].t_rxd1[0][1] = 1269ns;
slave_timing[0][22].t_rxd1[1][0] = 1142ns;
slave_timing[0][22].t_rxd1[0][2] = 906ns;
slave_timing[0][22].t_rxd1[2][0] = 1436ns;
slave_timing[0][22].t_rxd2[0][2] = 1376ns;
slave_timing[0][22].t_rxd2[2][0] = 948ns;
slave_timing[0][22].t_rxd2[1][2] = 1083ns;
slave_timing[0][22].t_rxd2[2][1] = 1363ns;

slave_timing[0][23].info_corner          = 0;
slave_timing[0][23].info_temp__j__       = 25;
slave_timing[0][23].info_i__quite_rec__  = 0.003000000;
slave_timing[0][23].info_dtr__ib__       = 1;
slave_timing[0][23].info_i__offset_rec__ = 0.001000000;
slave_timing[0][23].info_i__max_slave__  = 0.027000000;
slave_timing[0][23].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][23].info_r__dsi_bus__    = 5.000;

slave_timing[0][23].t_rxd1[0][1] = 1114ns;
slave_timing[0][23].t_rxd1[1][0] = 1303ns;
slave_timing[0][23].t_rxd1[0][2] = 834ns;
slave_timing[0][23].t_rxd1[2][0] = 1576ns;
slave_timing[0][23].t_rxd2[0][2] = 1270ns;
slave_timing[0][23].t_rxd2[2][0] = 1009ns;
slave_timing[0][23].t_rxd2[1][2] = 953ns;
slave_timing[0][23].t_rxd2[2][1] = 1640ns;

slave_timing[0][24].info_corner          = 0;
slave_timing[0][24].info_temp__j__       = 25;
slave_timing[0][24].info_i__quite_rec__  = 0.003000000;
slave_timing[0][24].info_dtr__ib__       = -1;
slave_timing[0][24].info_i__offset_rec__ = -0.001000000;
slave_timing[0][24].info_i__max_slave__  = 0.021000000;
slave_timing[0][24].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][24].info_r__dsi_bus__    = 5.000;

slave_timing[0][24].t_rxd1[0][1] = 1782ns;
slave_timing[0][24].t_rxd1[1][0] = 1249ns;
slave_timing[0][24].t_rxd1[0][2] = 1179ns;
slave_timing[0][24].t_rxd1[2][0] = 1605ns;
slave_timing[0][24].t_rxd2[0][2] = 2135ns;
slave_timing[0][24].t_rxd2[2][0] = 963ns;
slave_timing[0][24].t_rxd2[1][2] = 1805ns;
slave_timing[0][24].t_rxd2[2][1] = 1254ns;

slave_timing[0][25].info_corner          = 0;
slave_timing[0][25].info_temp__j__       = 25;
slave_timing[0][25].info_i__quite_rec__  = 0.003000000;
slave_timing[0][25].info_dtr__ib__       = -1;
slave_timing[0][25].info_i__offset_rec__ = 0.001000000;
slave_timing[0][25].info_i__max_slave__  = 0.021000000;
slave_timing[0][25].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][25].info_r__dsi_bus__    = 5.000;

slave_timing[0][25].t_rxd1[0][1] = 1450ns;
slave_timing[0][25].t_rxd1[1][0] = 1499ns;
slave_timing[0][25].t_rxd1[0][2] = 1058ns;
slave_timing[0][25].t_rxd1[2][0] = 1829ns;
slave_timing[0][25].t_rxd2[0][2] = 1784ns;
slave_timing[0][25].t_rxd2[2][0] = 1089ns;
slave_timing[0][25].t_rxd2[1][2] = 1461ns;
slave_timing[0][25].t_rxd2[2][1] = 1505ns;

slave_timing[0][26].info_corner          = 0;
slave_timing[0][26].info_temp__j__       = 25;
slave_timing[0][26].info_i__quite_rec__  = 0.003000000;
slave_timing[0][26].info_dtr__ib__       = -1;
slave_timing[0][26].info_i__offset_rec__ = -0.001000000;
slave_timing[0][26].info_i__max_slave__  = 0.027000000;
slave_timing[0][26].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][26].info_r__dsi_bus__    = 5.000;

slave_timing[0][26].t_rxd1[0][1] = 1460ns;
slave_timing[0][26].t_rxd1[1][0] = 1391ns;
slave_timing[0][26].t_rxd1[0][2] = 1063ns;
slave_timing[0][26].t_rxd1[2][0] = 1738ns;
slave_timing[0][26].t_rxd2[0][2] = 1569ns;
slave_timing[0][26].t_rxd2[2][0] = 1171ns;
slave_timing[0][26].t_rxd2[1][2] = 1188ns;
slave_timing[0][26].t_rxd2[2][1] = 1780ns;

slave_timing[0][27].info_corner          = 0;
slave_timing[0][27].info_temp__j__       = 25;
slave_timing[0][27].info_i__quite_rec__  = 0.003000000;
slave_timing[0][27].info_dtr__ib__       = -1;
slave_timing[0][27].info_i__offset_rec__ = 0.001000000;
slave_timing[0][27].info_i__max_slave__  = 0.027000000;
slave_timing[0][27].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][27].info_r__dsi_bus__    = 5.000;

slave_timing[0][27].t_rxd1[0][1] = 1271ns;
slave_timing[0][27].t_rxd1[1][0] = 1621ns;
slave_timing[0][27].t_rxd1[0][2] = 975ns;
slave_timing[0][27].t_rxd1[2][0] = 1936ns;
slave_timing[0][27].t_rxd2[0][2] = 1454ns;
slave_timing[0][27].t_rxd2[2][0] = 1257ns;
slave_timing[0][27].t_rxd2[1][2] = 1016ns;
slave_timing[0][27].t_rxd2[2][1] = 2387ns;

slave_timing[0][28].info_corner          = 0;
slave_timing[0][28].info_temp__j__       = 25;
slave_timing[0][28].info_i__quite_rec__  = 0.003000000;
slave_timing[0][28].info_dtr__ib__       = 1;
slave_timing[0][28].info_i__offset_rec__ = -0.001000000;
slave_timing[0][28].info_i__max_slave__  = 0.021000000;
slave_timing[0][28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][28].info_r__dsi_bus__    = 5.000;

slave_timing[0][28].t_rxd1[0][1] = 1899ns;
slave_timing[0][28].t_rxd1[1][0] = 1215ns;
slave_timing[0][28].t_rxd1[0][2] = 1196ns;
slave_timing[0][28].t_rxd1[2][0] = 1596ns;
slave_timing[0][28].t_rxd2[0][2] = 2450ns;
slave_timing[0][28].t_rxd2[2][0] = 915ns;
slave_timing[0][28].t_rxd2[1][2] = 2181ns;
slave_timing[0][28].t_rxd2[2][1] = 1145ns;

slave_timing[0][29].info_corner          = 0;
slave_timing[0][29].info_temp__j__       = 25;
slave_timing[0][29].info_i__quite_rec__  = 0.003000000;
slave_timing[0][29].info_dtr__ib__       = 1;
slave_timing[0][29].info_i__offset_rec__ = 0.001000000;
slave_timing[0][29].info_i__max_slave__  = 0.021000000;
slave_timing[0][29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][29].info_r__dsi_bus__    = 5.000;

slave_timing[0][29].t_rxd1[0][1] = 1515ns;
slave_timing[0][29].t_rxd1[1][0] = 1457ns;
slave_timing[0][29].t_rxd1[0][2] = 1085ns;
slave_timing[0][29].t_rxd1[2][0] = 1793ns;
slave_timing[0][29].t_rxd2[0][2] = 1940ns;
slave_timing[0][29].t_rxd2[2][0] = 1034ns;
slave_timing[0][29].t_rxd2[1][2] = 1640ns;
slave_timing[0][29].t_rxd2[2][1] = 1373ns;

slave_timing[0][30].info_corner          = 0;
slave_timing[0][30].info_temp__j__       = 25;
slave_timing[0][30].info_i__quite_rec__  = 0.003000000;
slave_timing[0][30].info_dtr__ib__       = 1;
slave_timing[0][30].info_i__offset_rec__ = -0.001000000;
slave_timing[0][30].info_i__max_slave__  = 0.027000000;
slave_timing[0][30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][30].info_r__dsi_bus__    = 5.000;

slave_timing[0][30].t_rxd1[0][1] = 1513ns;
slave_timing[0][30].t_rxd1[1][0] = 1364ns;
slave_timing[0][30].t_rxd1[0][2] = 1084ns;
slave_timing[0][30].t_rxd1[2][0] = 1714ns;
slave_timing[0][30].t_rxd2[0][2] = 1645ns;
slave_timing[0][30].t_rxd2[2][0] = 1130ns;
slave_timing[0][30].t_rxd2[1][2] = 1294ns;
slave_timing[0][30].t_rxd2[2][1] = 1631ns;

slave_timing[0][31].info_corner          = 0;
slave_timing[0][31].info_temp__j__       = 25;
slave_timing[0][31].info_i__quite_rec__  = 0.003000000;
slave_timing[0][31].info_dtr__ib__       = 1;
slave_timing[0][31].info_i__offset_rec__ = 0.001000000;
slave_timing[0][31].info_i__max_slave__  = 0.027000000;
slave_timing[0][31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][31].info_r__dsi_bus__    = 5.000;

slave_timing[0][31].t_rxd1[0][1] = 1331ns;
slave_timing[0][31].t_rxd1[1][0] = 1556ns;
slave_timing[0][31].t_rxd1[0][2] = 1006ns;
slave_timing[0][31].t_rxd1[2][0] = 1878ns;
slave_timing[0][31].t_rxd2[0][2] = 1529ns;
slave_timing[0][31].t_rxd2[2][0] = 1205ns;
slave_timing[0][31].t_rxd2[1][2] = 1137ns;
slave_timing[0][31].t_rxd2[2][1] = 1946ns;

slave_timing[0][32].info_corner          = 0;
slave_timing[0][32].info_temp__j__       = 25;
slave_timing[0][32].info_i__quite_rec__  = 0.000000000;
slave_timing[0][32].info_dtr__ib__       = -1;
slave_timing[0][32].info_i__offset_rec__ = -0.001000000;
slave_timing[0][32].info_i__max_slave__  = 0.021000000;
slave_timing[0][32].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][32].info_r__dsi_bus__    = 5.000;

slave_timing[0][32].t_rxd1[0][1] = 1519ns;
slave_timing[0][32].t_rxd1[1][0] = 1040ns;
slave_timing[0][32].t_rxd1[0][2] = 984ns;
slave_timing[0][32].t_rxd1[2][0] = 1352ns;
slave_timing[0][32].t_rxd2[0][2] = 1787ns;
slave_timing[0][32].t_rxd2[2][0] = 809ns;
slave_timing[0][32].t_rxd2[1][2] = 1534ns;
slave_timing[0][32].t_rxd2[2][1] = 1042ns;

slave_timing[0][33].info_corner          = 0;
slave_timing[0][33].info_temp__j__       = 25;
slave_timing[0][33].info_i__quite_rec__  = 0.000000000;
slave_timing[0][33].info_dtr__ib__       = -1;
slave_timing[0][33].info_i__offset_rec__ = 0.001000000;
slave_timing[0][33].info_i__max_slave__  = 0.021000000;
slave_timing[0][33].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][33].info_r__dsi_bus__    = 5.000;

slave_timing[0][33].t_rxd1[0][1] = 1225ns;
slave_timing[0][33].t_rxd1[1][0] = 1245ns;
slave_timing[0][33].t_rxd1[0][2] = 891ns;
slave_timing[0][33].t_rxd1[2][0] = 1528ns;
slave_timing[0][33].t_rxd2[0][2] = 1508ns;
slave_timing[0][33].t_rxd2[2][0] = 909ns;
slave_timing[0][33].t_rxd2[1][2] = 1239ns;
slave_timing[0][33].t_rxd2[2][1] = 1250ns;

slave_timing[0][34].info_corner          = 0;
slave_timing[0][34].info_temp__j__       = 25;
slave_timing[0][34].info_i__quite_rec__  = 0.000000000;
slave_timing[0][34].info_dtr__ib__       = -1;
slave_timing[0][34].info_i__offset_rec__ = -0.001000000;
slave_timing[0][34].info_i__max_slave__  = 0.027000000;
slave_timing[0][34].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][34].info_r__dsi_bus__    = 5.000;

slave_timing[0][34].t_rxd1[0][1] = 1234ns;
slave_timing[0][34].t_rxd1[1][0] = 1160ns;
slave_timing[0][34].t_rxd1[0][2] = 900ns;
slave_timing[0][34].t_rxd1[2][0] = 1450ns;
slave_timing[0][34].t_rxd2[0][2] = 1328ns;
slave_timing[0][34].t_rxd2[2][0] = 976ns;
slave_timing[0][34].t_rxd2[1][2] = 1007ns;
slave_timing[0][34].t_rxd2[2][1] = 1481ns;

slave_timing[0][35].info_corner          = 0;
slave_timing[0][35].info_temp__j__       = 25;
slave_timing[0][35].info_i__quite_rec__  = 0.000000000;
slave_timing[0][35].info_dtr__ib__       = -1;
slave_timing[0][35].info_i__offset_rec__ = 0.001000000;
slave_timing[0][35].info_i__max_slave__  = 0.027000000;
slave_timing[0][35].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][35].info_r__dsi_bus__    = 5.000;

slave_timing[0][35].t_rxd1[0][1] = 1069ns;
slave_timing[0][35].t_rxd1[1][0] = 1348ns;
slave_timing[0][35].t_rxd1[0][2] = 816ns;
slave_timing[0][35].t_rxd1[2][0] = 1622ns;
slave_timing[0][35].t_rxd2[0][2] = 1220ns;
slave_timing[0][35].t_rxd2[2][0] = 1050ns;
slave_timing[0][35].t_rxd2[1][2] = 861ns;
slave_timing[0][35].t_rxd2[2][1] = 1986ns;

slave_timing[0][36].info_corner          = 0;
slave_timing[0][36].info_temp__j__       = 25;
slave_timing[0][36].info_i__quite_rec__  = 0.000000000;
slave_timing[0][36].info_dtr__ib__       = 1;
slave_timing[0][36].info_i__offset_rec__ = -0.001000000;
slave_timing[0][36].info_i__max_slave__  = 0.021000000;
slave_timing[0][36].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][36].info_r__dsi_bus__    = 5.000;

slave_timing[0][36].t_rxd1[0][1] = 1687ns;
slave_timing[0][36].t_rxd1[1][0] = 992ns;
slave_timing[0][36].t_rxd1[0][2] = 1016ns;
slave_timing[0][36].t_rxd1[2][0] = 1316ns;
slave_timing[0][36].t_rxd2[0][2] = 2259ns;
slave_timing[0][36].t_rxd2[2][0] = 747ns;
slave_timing[0][36].t_rxd2[1][2] = 2021ns;
slave_timing[0][36].t_rxd2[2][1] = 932ns;

slave_timing[0][37].info_corner          = 0;
slave_timing[0][37].info_temp__j__       = 25;
slave_timing[0][37].info_i__quite_rec__  = 0.000000000;
slave_timing[0][37].info_dtr__ib__       = 1;
slave_timing[0][37].info_i__offset_rec__ = 0.001000000;
slave_timing[0][37].info_i__max_slave__  = 0.021000000;
slave_timing[0][37].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][37].info_r__dsi_bus__    = 5.000;

slave_timing[0][37].t_rxd1[0][1] = 1310ns;
slave_timing[0][37].t_rxd1[1][0] = 1186ns;
slave_timing[0][37].t_rxd1[0][2] = 924ns;
slave_timing[0][37].t_rxd1[2][0] = 1474ns;
slave_timing[0][37].t_rxd2[0][2] = 1681ns;
slave_timing[0][37].t_rxd2[2][0] = 851ns;
slave_timing[0][37].t_rxd2[1][2] = 1425ns;
slave_timing[0][37].t_rxd2[2][1] = 1120ns;

slave_timing[0][38].info_corner          = 0;
slave_timing[0][38].info_temp__j__       = 25;
slave_timing[0][38].info_i__quite_rec__  = 0.000000000;
slave_timing[0][38].info_dtr__ib__       = 1;
slave_timing[0][38].info_i__offset_rec__ = -0.001000000;
slave_timing[0][38].info_i__max_slave__  = 0.027000000;
slave_timing[0][38].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][38].info_r__dsi_bus__    = 5.000;

slave_timing[0][38].t_rxd1[0][1] = 1297ns;
slave_timing[0][38].t_rxd1[1][0] = 1117ns;
slave_timing[0][38].t_rxd1[0][2] = 919ns;
slave_timing[0][38].t_rxd1[2][0] = 1415ns;
slave_timing[0][38].t_rxd2[0][2] = 1399ns;
slave_timing[0][38].t_rxd2[2][0] = 934ns;
slave_timing[0][38].t_rxd2[1][2] = 1107ns;
slave_timing[0][38].t_rxd2[2][1] = 1329ns;

slave_timing[0][39].info_corner          = 0;
slave_timing[0][39].info_temp__j__       = 25;
slave_timing[0][39].info_i__quite_rec__  = 0.000000000;
slave_timing[0][39].info_dtr__ib__       = 1;
slave_timing[0][39].info_i__offset_rec__ = 0.001000000;
slave_timing[0][39].info_i__max_slave__  = 0.027000000;
slave_timing[0][39].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][39].info_r__dsi_bus__    = 5.000;

slave_timing[0][39].t_rxd1[0][1] = 1125ns;
slave_timing[0][39].t_rxd1[1][0] = 1291ns;
slave_timing[0][39].t_rxd1[0][2] = 844ns;
slave_timing[0][39].t_rxd1[2][0] = 1567ns;
slave_timing[0][39].t_rxd2[0][2] = 1286ns;
slave_timing[0][39].t_rxd2[2][0] = 1004ns;
slave_timing[0][39].t_rxd2[1][2] = 963ns;
slave_timing[0][39].t_rxd2[2][1] = 1616ns;

slave_timing[0][40].info_corner          = 0;
slave_timing[0][40].info_temp__j__       = 25;
slave_timing[0][40].info_i__quite_rec__  = 0.000000000;
slave_timing[0][40].info_dtr__ib__       = -1;
slave_timing[0][40].info_i__offset_rec__ = -0.001000000;
slave_timing[0][40].info_i__max_slave__  = 0.021000000;
slave_timing[0][40].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][40].info_r__dsi_bus__    = 5.000;

slave_timing[0][40].t_rxd1[0][1] = 1807ns;
slave_timing[0][40].t_rxd1[1][0] = 1240ns;
slave_timing[0][40].t_rxd1[0][2] = 1183ns;
slave_timing[0][40].t_rxd1[2][0] = 1617ns;
slave_timing[0][40].t_rxd2[0][2] = 2159ns;
slave_timing[0][40].t_rxd2[2][0] = 971ns;
slave_timing[0][40].t_rxd2[1][2] = 1827ns;
slave_timing[0][40].t_rxd2[2][1] = 1243ns;

slave_timing[0][41].info_corner          = 0;
slave_timing[0][41].info_temp__j__       = 25;
slave_timing[0][41].info_i__quite_rec__  = 0.000000000;
slave_timing[0][41].info_dtr__ib__       = -1;
slave_timing[0][41].info_i__offset_rec__ = 0.001000000;
slave_timing[0][41].info_i__max_slave__  = 0.021000000;
slave_timing[0][41].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][41].info_r__dsi_bus__    = 5.000;

slave_timing[0][41].t_rxd1[0][1] = 1462ns;
slave_timing[0][41].t_rxd1[1][0] = 1488ns;
slave_timing[0][41].t_rxd1[0][2] = 1065ns;
slave_timing[0][41].t_rxd1[2][0] = 1819ns;
slave_timing[0][41].t_rxd2[0][2] = 1798ns;
slave_timing[0][41].t_rxd2[2][0] = 1083ns;
slave_timing[0][41].t_rxd2[1][2] = 1475ns;
slave_timing[0][41].t_rxd2[2][1] = 1492ns;

slave_timing[0][42].info_corner          = 0;
slave_timing[0][42].info_temp__j__       = 25;
slave_timing[0][42].info_i__quite_rec__  = 0.000000000;
slave_timing[0][42].info_dtr__ib__       = -1;
slave_timing[0][42].info_i__offset_rec__ = -0.001000000;
slave_timing[0][42].info_i__max_slave__  = 0.027000000;
slave_timing[0][42].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][42].info_r__dsi_bus__    = 5.000;

slave_timing[0][42].t_rxd1[0][1] = 1473ns;
slave_timing[0][42].t_rxd1[1][0] = 1386ns;
slave_timing[0][42].t_rxd1[0][2] = 1074ns;
slave_timing[0][42].t_rxd1[2][0] = 1716ns;
slave_timing[0][42].t_rxd2[0][2] = 1588ns;
slave_timing[0][42].t_rxd2[2][0] = 1159ns;
slave_timing[0][42].t_rxd2[1][2] = 1199ns;
slave_timing[0][42].t_rxd2[2][1] = 1765ns;

slave_timing[0][43].info_corner          = 0;
slave_timing[0][43].info_temp__j__       = 25;
slave_timing[0][43].info_i__quite_rec__  = 0.000000000;
slave_timing[0][43].info_dtr__ib__       = -1;
slave_timing[0][43].info_i__offset_rec__ = 0.001000000;
slave_timing[0][43].info_i__max_slave__  = 0.027000000;
slave_timing[0][43].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][43].info_r__dsi_bus__    = 5.000;

slave_timing[0][43].t_rxd1[0][1] = 1279ns;
slave_timing[0][43].t_rxd1[1][0] = 1609ns;
slave_timing[0][43].t_rxd1[0][2] = 979ns;
slave_timing[0][43].t_rxd1[2][0] = 1928ns;
slave_timing[0][43].t_rxd2[0][2] = 1460ns;
slave_timing[0][43].t_rxd2[2][0] = 1253ns;
slave_timing[0][43].t_rxd2[1][2] = 1025ns;
slave_timing[0][43].t_rxd2[2][1] = 2333ns;

slave_timing[0][44].info_corner          = 0;
slave_timing[0][44].info_temp__j__       = 25;
slave_timing[0][44].info_i__quite_rec__  = 0.000000000;
slave_timing[0][44].info_dtr__ib__       = 1;
slave_timing[0][44].info_i__offset_rec__ = -0.001000000;
slave_timing[0][44].info_i__max_slave__  = 0.021000000;
slave_timing[0][44].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][44].info_r__dsi_bus__    = 5.000;

slave_timing[0][44].t_rxd1[0][1] = 1997ns;
slave_timing[0][44].t_rxd1[1][0] = 1183ns;
slave_timing[0][44].t_rxd1[0][2] = 1213ns;
slave_timing[0][44].t_rxd1[2][0] = 1571ns;
slave_timing[0][44].t_rxd2[0][2] = 2634ns;
slave_timing[0][44].t_rxd2[2][0] = 894ns;
slave_timing[0][44].t_rxd2[1][2] = 2374ns;
slave_timing[0][44].t_rxd2[2][1] = 1111ns;

slave_timing[0][45].info_corner          = 0;
slave_timing[0][45].info_temp__j__       = 25;
slave_timing[0][45].info_i__quite_rec__  = 0.000000000;
slave_timing[0][45].info_dtr__ib__       = 1;
slave_timing[0][45].info_i__offset_rec__ = 0.001000000;
slave_timing[0][45].info_i__max_slave__  = 0.021000000;
slave_timing[0][45].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][45].info_r__dsi_bus__    = 5.000;

slave_timing[0][45].t_rxd1[0][1] = 1562ns;
slave_timing[0][45].t_rxd1[1][0] = 1414ns;
slave_timing[0][45].t_rxd1[0][2] = 1102ns;
slave_timing[0][45].t_rxd1[2][0] = 1758ns;
slave_timing[0][45].t_rxd2[0][2] = 1993ns;
slave_timing[0][45].t_rxd2[2][0] = 1018ns;
slave_timing[0][45].t_rxd2[1][2] = 1698ns;
slave_timing[0][45].t_rxd2[2][1] = 1337ns;

slave_timing[0][46].info_corner          = 0;
slave_timing[0][46].info_temp__j__       = 25;
slave_timing[0][46].info_i__quite_rec__  = 0.000000000;
slave_timing[0][46].info_dtr__ib__       = 1;
slave_timing[0][46].info_i__offset_rec__ = -0.001000000;
slave_timing[0][46].info_i__max_slave__  = 0.027000000;
slave_timing[0][46].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][46].info_r__dsi_bus__    = 5.000;

slave_timing[0][46].t_rxd1[0][1] = 1527ns;
slave_timing[0][46].t_rxd1[1][0] = 1355ns;
slave_timing[0][46].t_rxd1[0][2] = 1089ns;
slave_timing[0][46].t_rxd1[2][0] = 1707ns;
slave_timing[0][46].t_rxd2[0][2] = 1656ns;
slave_timing[0][46].t_rxd2[2][0] = 1124ns;
slave_timing[0][46].t_rxd2[1][2] = 1303ns;
slave_timing[0][46].t_rxd2[2][1] = 1612ns;

slave_timing[0][47].info_corner          = 0;
slave_timing[0][47].info_temp__j__       = 25;
slave_timing[0][47].info_i__quite_rec__  = 0.000000000;
slave_timing[0][47].info_dtr__ib__       = 1;
slave_timing[0][47].info_i__offset_rec__ = 0.001000000;
slave_timing[0][47].info_i__max_slave__  = 0.027000000;
slave_timing[0][47].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][47].info_r__dsi_bus__    = 5.000;

slave_timing[0][47].t_rxd1[0][1] = 1323ns;
slave_timing[0][47].t_rxd1[1][0] = 1570ns;
slave_timing[0][47].t_rxd1[0][2] = 999ns;
slave_timing[0][47].t_rxd1[2][0] = 1891ns;
slave_timing[0][47].t_rxd2[0][2] = 1524ns;
slave_timing[0][47].t_rxd2[2][0] = 1209ns;
slave_timing[0][47].t_rxd2[1][2] = 1132ns;
slave_timing[0][47].t_rxd2[2][1] = 1970ns;

slave_timing[0][48].info_corner          = 0;
slave_timing[0][48].info_temp__j__       = 25;
slave_timing[0][48].info_i__quite_rec__  = 0.040000000;
slave_timing[0][48].info_dtr__ib__       = -1;
slave_timing[0][48].info_i__offset_rec__ = -0.001000000;
slave_timing[0][48].info_i__max_slave__  = 0.021000000;
slave_timing[0][48].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][48].info_r__dsi_bus__    = 5.000;

slave_timing[0][48].t_rxd1[0][1] = 1406ns;
slave_timing[0][48].t_rxd1[1][0] = 1101ns;
slave_timing[0][48].t_rxd1[0][2] = 955ns;
slave_timing[0][48].t_rxd1[2][0] = 1400ns;
slave_timing[0][48].t_rxd2[0][2] = 1676ns;
slave_timing[0][48].t_rxd2[2][0] = 842ns;
slave_timing[0][48].t_rxd2[1][2] = 1421ns;
slave_timing[0][48].t_rxd2[2][1] = 1102ns;

slave_timing[0][49].info_corner          = 0;
slave_timing[0][49].info_temp__j__       = 25;
slave_timing[0][49].info_i__quite_rec__  = 0.040000000;
slave_timing[0][49].info_dtr__ib__       = -1;
slave_timing[0][49].info_i__offset_rec__ = 0.001000000;
slave_timing[0][49].info_i__max_slave__  = 0.021000000;
slave_timing[0][49].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][49].info_r__dsi_bus__    = 5.000;

slave_timing[0][49].t_rxd1[0][1] = 1157ns;
slave_timing[0][49].t_rxd1[1][0] = 1326ns;
slave_timing[0][49].t_rxd1[0][2] = 862ns;
slave_timing[0][49].t_rxd1[2][0] = 1597ns;
slave_timing[0][49].t_rxd2[0][2] = 1447ns;
slave_timing[0][49].t_rxd2[2][0] = 935ns;
slave_timing[0][49].t_rxd2[1][2] = 1166ns;
slave_timing[0][49].t_rxd2[2][1] = 1327ns;

slave_timing[0][50].info_corner          = 0;
slave_timing[0][50].info_temp__j__       = 25;
slave_timing[0][50].info_i__quite_rec__  = 0.040000000;
slave_timing[0][50].info_dtr__ib__       = -1;
slave_timing[0][50].info_i__offset_rec__ = -0.001000000;
slave_timing[0][50].info_i__max_slave__  = 0.027000000;
slave_timing[0][50].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][50].info_r__dsi_bus__    = 5.000;

slave_timing[0][50].t_rxd1[0][1] = 1212ns;
slave_timing[0][50].t_rxd1[1][0] = 1183ns;
slave_timing[0][50].t_rxd1[0][2] = 885ns;
slave_timing[0][50].t_rxd1[2][0] = 1469ns;
slave_timing[0][50].t_rxd2[0][2] = 1305ns;
slave_timing[0][50].t_rxd2[2][0] = 986ns;
slave_timing[0][50].t_rxd2[1][2] = 987ns;
slave_timing[0][50].t_rxd2[2][1] = 1515ns;

slave_timing[0][51].info_corner          = 0;
slave_timing[0][51].info_temp__j__       = 25;
slave_timing[0][51].info_i__quite_rec__  = 0.040000000;
slave_timing[0][51].info_dtr__ib__       = -1;
slave_timing[0][51].info_i__offset_rec__ = 0.001000000;
slave_timing[0][51].info_i__max_slave__  = 0.027000000;
slave_timing[0][51].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][51].info_r__dsi_bus__    = 5.000;

slave_timing[0][51].t_rxd1[0][1] = 1069ns;
slave_timing[0][51].t_rxd1[1][0] = 1358ns;
slave_timing[0][51].t_rxd1[0][2] = 808ns;
slave_timing[0][51].t_rxd1[2][0] = 1627ns;
slave_timing[0][51].t_rxd2[0][2] = 1209ns;
slave_timing[0][51].t_rxd2[2][0] = 1049ns;
slave_timing[0][51].t_rxd2[1][2] = 856ns;
slave_timing[0][51].t_rxd2[2][1] = 2002ns;

slave_timing[0][52].info_corner          = 0;
slave_timing[0][52].info_temp__j__       = 25;
slave_timing[0][52].info_i__quite_rec__  = 0.040000000;
slave_timing[0][52].info_dtr__ib__       = 1;
slave_timing[0][52].info_i__offset_rec__ = -0.001000000;
slave_timing[0][52].info_i__max_slave__  = 0.021000000;
slave_timing[0][52].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][52].info_r__dsi_bus__    = 5.000;

slave_timing[0][52].t_rxd1[0][1] = 1645ns;
slave_timing[0][52].t_rxd1[1][0] = 1005ns;
slave_timing[0][52].t_rxd1[0][2] = 1010ns;
slave_timing[0][52].t_rxd1[2][0] = 1325ns;
slave_timing[0][52].t_rxd2[0][2] = 2174ns;
slave_timing[0][52].t_rxd2[2][0] = 756ns;
slave_timing[0][52].t_rxd2[1][2] = 1935ns;
slave_timing[0][52].t_rxd2[2][1] = 948ns;

slave_timing[0][53].info_corner          = 0;
slave_timing[0][53].info_temp__j__       = 25;
slave_timing[0][53].info_i__quite_rec__  = 0.040000000;
slave_timing[0][53].info_dtr__ib__       = 1;
slave_timing[0][53].info_i__offset_rec__ = 0.001000000;
slave_timing[0][53].info_i__max_slave__  = 0.021000000;
slave_timing[0][53].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][53].info_r__dsi_bus__    = 5.000;

slave_timing[0][53].t_rxd1[0][1] = 1291ns;
slave_timing[0][53].t_rxd1[1][0] = 1201ns;
slave_timing[0][53].t_rxd1[0][2] = 917ns;
slave_timing[0][53].t_rxd1[2][0] = 1488ns;
slave_timing[0][53].t_rxd2[0][2] = 1657ns;
slave_timing[0][53].t_rxd2[2][0] = 860ns;
slave_timing[0][53].t_rxd2[1][2] = 1400ns;
slave_timing[0][53].t_rxd2[2][1] = 1133ns;

slave_timing[0][54].info_corner          = 0;
slave_timing[0][54].info_temp__j__       = 25;
slave_timing[0][54].info_i__quite_rec__  = 0.040000000;
slave_timing[0][54].info_dtr__ib__       = 1;
slave_timing[0][54].info_i__offset_rec__ = -0.001000000;
slave_timing[0][54].info_i__max_slave__  = 0.027000000;
slave_timing[0][54].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][54].info_r__dsi_bus__    = 5.000;

slave_timing[0][54].t_rxd1[0][1] = 1306ns;
slave_timing[0][54].t_rxd1[1][0] = 1112ns;
slave_timing[0][54].t_rxd1[0][2] = 921ns;
slave_timing[0][54].t_rxd1[2][0] = 1411ns;
slave_timing[0][54].t_rxd2[0][2] = 1401ns;
slave_timing[0][54].t_rxd2[2][0] = 934ns;
slave_timing[0][54].t_rxd2[1][2] = 1113ns;
slave_timing[0][54].t_rxd2[2][1] = 1322ns;

slave_timing[0][55].info_corner          = 0;
slave_timing[0][55].info_temp__j__       = 25;
slave_timing[0][55].info_i__quite_rec__  = 0.040000000;
slave_timing[0][55].info_dtr__ib__       = 1;
slave_timing[0][55].info_i__offset_rec__ = 0.001000000;
slave_timing[0][55].info_i__max_slave__  = 0.027000000;
slave_timing[0][55].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][55].info_r__dsi_bus__    = 5.000;

slave_timing[0][55].t_rxd1[0][1] = 1130ns;
slave_timing[0][55].t_rxd1[1][0] = 1285ns;
slave_timing[0][55].t_rxd1[0][2] = 847ns;
slave_timing[0][55].t_rxd1[2][0] = 1563ns;
slave_timing[0][55].t_rxd2[0][2] = 1288ns;
slave_timing[0][55].t_rxd2[2][0] = 1005ns;
slave_timing[0][55].t_rxd2[1][2] = 965ns;
slave_timing[0][55].t_rxd2[2][1] = 1604ns;

slave_timing[0][56].info_corner          = 0;
slave_timing[0][56].info_temp__j__       = 25;
slave_timing[0][56].info_i__quite_rec__  = 0.040000000;
slave_timing[0][56].info_dtr__ib__       = -1;
slave_timing[0][56].info_i__offset_rec__ = -0.001000000;
slave_timing[0][56].info_i__max_slave__  = 0.021000000;
slave_timing[0][56].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][56].info_r__dsi_bus__    = 5.000;

slave_timing[0][56].t_rxd1[0][1] = 1675ns;
slave_timing[0][56].t_rxd1[1][0] = 1313ns;
slave_timing[0][56].t_rxd1[0][2] = 1139ns;
slave_timing[0][56].t_rxd1[2][0] = 1673ns;
slave_timing[0][56].t_rxd2[0][2] = 1991ns;
slave_timing[0][56].t_rxd2[2][0] = 1007ns;
slave_timing[0][56].t_rxd2[1][2] = 1693ns;
slave_timing[0][56].t_rxd2[2][1] = 1316ns;

slave_timing[0][57].info_corner          = 0;
slave_timing[0][57].info_temp__j__       = 25;
slave_timing[0][57].info_i__quite_rec__  = 0.040000000;
slave_timing[0][57].info_dtr__ib__       = -1;
slave_timing[0][57].info_i__offset_rec__ = 0.001000000;
slave_timing[0][57].info_i__max_slave__  = 0.021000000;
slave_timing[0][57].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][57].info_r__dsi_bus__    = 5.000;

slave_timing[0][57].t_rxd1[0][1] = 1377ns;
slave_timing[0][57].t_rxd1[1][0] = 1583ns;
slave_timing[0][57].t_rxd1[0][2] = 1028ns;
slave_timing[0][57].t_rxd1[2][0] = 1905ns;
slave_timing[0][57].t_rxd2[0][2] = 1726ns;
slave_timing[0][57].t_rxd2[2][0] = 1119ns;
slave_timing[0][57].t_rxd2[1][2] = 1390ns;
slave_timing[0][57].t_rxd2[2][1] = 1586ns;

slave_timing[0][58].info_corner          = 0;
slave_timing[0][58].info_temp__j__       = 25;
slave_timing[0][58].info_i__quite_rec__  = 0.040000000;
slave_timing[0][58].info_dtr__ib__       = -1;
slave_timing[0][58].info_i__offset_rec__ = -0.001000000;
slave_timing[0][58].info_i__max_slave__  = 0.027000000;
slave_timing[0][58].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][58].info_r__dsi_bus__    = 5.000;

slave_timing[0][58].t_rxd1[0][1] = 1444ns;
slave_timing[0][58].t_rxd1[1][0] = 1414ns;
slave_timing[0][58].t_rxd1[0][2] = 1056ns;
slave_timing[0][58].t_rxd1[2][0] = 1755ns;
slave_timing[0][58].t_rxd2[0][2] = 1560ns;
slave_timing[0][58].t_rxd2[2][0] = 1178ns;
slave_timing[0][58].t_rxd2[1][2] = 1179ns;
slave_timing[0][58].t_rxd2[2][1] = 1808ns;

slave_timing[0][59].info_corner          = 0;
slave_timing[0][59].info_temp__j__       = 25;
slave_timing[0][59].info_i__quite_rec__  = 0.040000000;
slave_timing[0][59].info_dtr__ib__       = -1;
slave_timing[0][59].info_i__offset_rec__ = 0.001000000;
slave_timing[0][59].info_i__max_slave__  = 0.027000000;
slave_timing[0][59].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][59].info_r__dsi_bus__    = 5.000;

slave_timing[0][59].t_rxd1[0][1] = 1274ns;
slave_timing[0][59].t_rxd1[1][0] = 1622ns;
slave_timing[0][59].t_rxd1[0][2] = 964ns;
slave_timing[0][59].t_rxd1[2][0] = 1937ns;
slave_timing[0][59].t_rxd2[0][2] = 1444ns;
slave_timing[0][59].t_rxd2[2][0] = 1254ns;
slave_timing[0][59].t_rxd2[1][2] = 1021ns;
slave_timing[0][59].t_rxd2[2][1] = 2354ns;

slave_timing[0][60].info_corner          = 0;
slave_timing[0][60].info_temp__j__       = 25;
slave_timing[0][60].info_i__quite_rec__  = 0.040000000;
slave_timing[0][60].info_dtr__ib__       = 1;
slave_timing[0][60].info_i__offset_rec__ = -0.001000000;
slave_timing[0][60].info_i__max_slave__  = 0.021000000;
slave_timing[0][60].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][60].info_r__dsi_bus__    = 5.000;

slave_timing[0][60].t_rxd1[0][1] = 1950ns;
slave_timing[0][60].t_rxd1[1][0] = 1198ns;
slave_timing[0][60].t_rxd1[0][2] = 1207ns;
slave_timing[0][60].t_rxd1[2][0] = 1585ns;
slave_timing[0][60].t_rxd2[0][2] = 2543ns;
slave_timing[0][60].t_rxd2[2][0] = 906ns;
slave_timing[0][60].t_rxd2[1][2] = 2278ns;
slave_timing[0][60].t_rxd2[2][1] = 1127ns;

slave_timing[0][61].info_corner          = 0;
slave_timing[0][61].info_temp__j__       = 25;
slave_timing[0][61].info_i__quite_rec__  = 0.040000000;
slave_timing[0][61].info_dtr__ib__       = 1;
slave_timing[0][61].info_i__offset_rec__ = 0.001000000;
slave_timing[0][61].info_i__max_slave__  = 0.021000000;
slave_timing[0][61].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][61].info_r__dsi_bus__    = 5.000;

slave_timing[0][61].t_rxd1[0][1] = 1541ns;
slave_timing[0][61].t_rxd1[1][0] = 1435ns;
slave_timing[0][61].t_rxd1[0][2] = 1096ns;
slave_timing[0][61].t_rxd1[2][0] = 1775ns;
slave_timing[0][61].t_rxd2[0][2] = 1972ns;
slave_timing[0][61].t_rxd2[2][0] = 1027ns;
slave_timing[0][61].t_rxd2[1][2] = 1670ns;
slave_timing[0][61].t_rxd2[2][1] = 1352ns;

slave_timing[0][62].info_corner          = 0;
slave_timing[0][62].info_temp__j__       = 25;
slave_timing[0][62].info_i__quite_rec__  = 0.040000000;
slave_timing[0][62].info_dtr__ib__       = 1;
slave_timing[0][62].info_i__offset_rec__ = -0.001000000;
slave_timing[0][62].info_i__max_slave__  = 0.027000000;
slave_timing[0][62].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][62].info_r__dsi_bus__    = 5.000;

slave_timing[0][62].t_rxd1[0][1] = 1558ns;
slave_timing[0][62].t_rxd1[1][0] = 1329ns;
slave_timing[0][62].t_rxd1[0][2] = 1101ns;
slave_timing[0][62].t_rxd1[2][0] = 1685ns;
slave_timing[0][62].t_rxd2[0][2] = 1675ns;
slave_timing[0][62].t_rxd2[2][0] = 1114ns;
slave_timing[0][62].t_rxd2[1][2] = 1327ns;
slave_timing[0][62].t_rxd2[2][1] = 1580ns;

slave_timing[0][63].info_corner          = 0;
slave_timing[0][63].info_temp__j__       = 25;
slave_timing[0][63].info_i__quite_rec__  = 0.040000000;
slave_timing[0][63].info_dtr__ib__       = 1;
slave_timing[0][63].info_i__offset_rec__ = 0.001000000;
slave_timing[0][63].info_i__max_slave__  = 0.027000000;
slave_timing[0][63].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][63].info_r__dsi_bus__    = 5.000;

slave_timing[0][63].t_rxd1[0][1] = 1351ns;
slave_timing[0][63].t_rxd1[1][0] = 1535ns;
slave_timing[0][63].t_rxd1[0][2] = 1013ns;
slave_timing[0][63].t_rxd1[2][0] = 1861ns;
slave_timing[0][63].t_rxd2[0][2] = 1539ns;
slave_timing[0][63].t_rxd2[2][0] = 1199ns;
slave_timing[0][63].t_rxd2[1][2] = 1153ns;
slave_timing[0][63].t_rxd2[2][1] = 1907ns;

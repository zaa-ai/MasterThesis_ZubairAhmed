/* ###   interface instances   ###################################################### */

OTP_readout_register_OTP_READ_ADDRESS_if OTP_readout_register_OTP_READ_ADDRESS (); 
OTP_readout_register_OTP_READ_VALUE_if OTP_readout_register_OTP_READ_VALUE (); 
OTP_readout_register_OTP_READ_STATUS_if OTP_readout_register_OTP_READ_STATUS (); 


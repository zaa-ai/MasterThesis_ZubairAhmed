task send_p52143_413_response();
	#	0us;	slave_if.cable.Current = 	0	;
	#	34.08us;	slave_if.cable.Current = 	1	;
	#	0.992us;	slave_if.cable.Current = 	2	;
	#	2.288us;	slave_if.cable.Current = 	1	;
	#	8.944us;	slave_if.cable.Current = 	0	;
	#	2.664us;	slave_if.cable.Current = 	1	;
	#	1.048us;	slave_if.cable.Current = 	2	;
	#	2.232us;	slave_if.cable.Current = 	1	;
	#	5.944us;	slave_if.cable.Current = 	0	;
	#	3.384us;	slave_if.cable.Current = 	1	;
	#	2.616us;	slave_if.cable.Current = 	0	;
	#	2.72us;	slave_if.cable.Current = 	1	;
	#	1.056us;	slave_if.cable.Current = 	2	;
	#	2.168us;	slave_if.cable.Current = 	1	;
	#	6us;	slave_if.cable.Current = 	0	;
	#	2.72us;	slave_if.cable.Current = 	1	;
	#	1us;	slave_if.cable.Current = 	2	;
	#	1.728us;	slave_if.cable.Current = 	1	;
	#	1.056us;	slave_if.cable.Current = 	0	;
	#	2.16us;	slave_if.cable.Current = 	1	;
	#	1.056us;	slave_if.cable.Current = 	2	;
	#	2.168us;	slave_if.cable.Current = 	1	;
	#	6us;	slave_if.cable.Current = 	0	;
	#	3.328us;	slave_if.cable.Current = 	1	;
	#	2.672us;	slave_if.cable.Current = 	0	;
	#	6.328us;	slave_if.cable.Current = 	1	;
	#	5.616us;	slave_if.cable.Current = 	0	;
	#	2.72us;	slave_if.cable.Current = 	1	;
	#	1.056us;	slave_if.cable.Current = 	2	;
	#	2.168us;	slave_if.cable.Current = 	1	;
	#	3.328us;	slave_if.cable.Current = 	2	;
	#	2.616us;	slave_if.cable.Current = 	1	;
	#	6.008us;	slave_if.cable.Current = 	0	;
	#	3.32us;	slave_if.cable.Current = 	1	;
	#	6us;	slave_if.cable.Current = 	2	;
	#	2.56us;	slave_if.cable.Current = 	1	;
	#	6.008us;	slave_if.cable.Current = 	0	;
	#	2.656us;	slave_if.cable.Current = 	1	;
	#	1.056us;	slave_if.cable.Current = 	2	;
	#	1.728us;	slave_if.cable.Current = 	1	;
	#	1us;	slave_if.cable.Current = 	0	;
	#	2.824us;	slave_if.cable.Current = 	1	;
	#	8.624us;	slave_if.cable.Current = 	0	;
	#	2.656us;	slave_if.cable.Current = 	1	;
	#	1.056us;	slave_if.cable.Current = 	2	;
	#	4.728us;	slave_if.cable.Current = 	1	;
	#	1us;	slave_if.cable.Current = 	0	;
	#	2.832us;	slave_if.cable.Current = 	1	;
	#	5.616us;	slave_if.cable.Current = 	0	;
	#	2.712us;	slave_if.cable.Current = 	1	;
	#	1.056us;	slave_if.cable.Current = 	2	;
	#	2.176us;	slave_if.cable.Current = 	1	;
	#	3us;	slave_if.cable.Current = 	0	;
	#	3.328us;	slave_if.cable.Current = 	1	;
	#	5.616us;	slave_if.cable.Current = 	0	;
	#	3.384us;	slave_if.cable.Current = 	1	;
	#	2.944us;	slave_if.cable.Current = 	2	;
	#	5.56us;	slave_if.cable.Current = 	1	;
	#	6us;	slave_if.cable.Current = 	0	;
	#	2.72us;	slave_if.cable.Current = 	1	;
	#	1us;	slave_if.cable.Current = 	2	;
	#	5.168us;	slave_if.cable.Current = 	1	;
	#	8.896us;	slave_if.cable.Current = 	0	;
	#	3.544us;	slave_if.cable.Current = 	1	;
	#	3us;	slave_if.cable.Current = 	2	;
	#	1.952us;	slave_if.cable.Current = 	1	;
	#	1us;	slave_if.cable.Current = 	0	;
	#	2.992us;	slave_if.cable.Current = 	1	;
	#	5.456us;	slave_if.cable.Current = 	0	;
	#	2.824us;	slave_if.cable.Current = 	1	;
	#	1.056us;	slave_if.cable.Current = 	2	;
	#	1.616us;	slave_if.cable.Current = 	1	;
	#	1us;	slave_if.cable.Current = 	0	;
	#	5.992us;	slave_if.cable.Current = 	1	;
	#	5.392us;	slave_if.cable.Current = 	0	;
	#	3.552us;	slave_if.cable.Current = 	1	;
	#	2.448us;	slave_if.cable.Current = 	0	;
	#	3.552us;	slave_if.cable.Current = 	1	;
	#	8.4us;	slave_if.cable.Current = 	0	;
	#	3.544us;	slave_if.cable.Current = 	1	;
	#	2.944us;	slave_if.cable.Current = 	2	;
	#	2.4us;	slave_if.cable.Current = 	1	;
	#	3.544us;	slave_if.cable.Current = 	2	;
	#	2.456us;	slave_if.cable.Current = 	1	;
	#	11.94399us;	slave_if.cable.Current = 	0	;
	#	2.824us;	slave_if.cable.Current = 	1	;
	#	1.056us;	slave_if.cable.Current = 	2	;
	#	2.064us;	slave_if.cable.Current = 	1	;
	#	6.488us;	slave_if.cable.Current = 	2	;
	#	2.4us;	slave_if.cable.Current = 	1	;
	#	6.544us;	slave_if.cable.Current = 	2	;
	#	2.4us;	slave_if.cable.Current = 	1	;
	#	8.944us;	slave_if.cable.Current = 	0	;
	#	2.88us;	slave_if.cable.Current = 	1	;
	#	1.056us;	slave_if.cable.Current = 	2	;
	#	4.952us;	slave_if.cable.Current = 	1	;
	#	6.552us;	slave_if.cable.Current = 	2	;
	#	1.952us;	slave_if.cable.Current = 	1	;
	#	1.056us;	slave_if.cable.Current = 	0	;
	#	2.272us;	slave_if.cable.Current = 	1	;
	#	1.056us;	slave_if.cable.Current = 	2	;
	#	4.888us;	slave_if.cable.Current = 	1	;
	#	9us;	slave_if.cable.Current = 	0	;
	#	5.936us;	slave_if.cable.Current = 	1	;
	#	1.112us;	slave_if.cable.Current = 	2	;
	#	1.84us;	slave_if.cable.Current = 	1	;
	#	6.832us;	slave_if.cable.Current = 	2	;
	#	2.12us;	slave_if.cable.Current = 	1	;
	#	3.768us;	slave_if.cable.Current = 	2	;
	#	5.12us;	slave_if.cable.Current = 	1	;
	#	12.768us;	slave_if.cable.Current = 	2	;
	#	5.12us;	slave_if.cable.Current = 	1	;
	#	6.712us;	slave_if.cable.Current = 	2	;
	#	1.784us;	slave_if.cable.Current = 	1	;
	#	1us;	slave_if.cable.Current = 	0	;
	#	3.216us;	slave_if.cable.Current = 	1	;
	#	3us;	slave_if.cable.Current = 	2	;
	#	2.176us;	slave_if.cable.Current = 	1	;
	#	6.712us;	slave_if.cable.Current = 	2	;
	#	4.728us;	slave_if.cable.Current = 	1	;
	#	1.056us;	slave_if.cable.Current = 	0	;
	#	2.328us;	slave_if.cable.Current = 	1	;
	#	1.168us;	slave_if.cable.Current = 	2	;
	#	1.84us;	slave_if.cable.Current = 	1	;
	#	6.768us;	slave_if.cable.Current = 	2	;
	#	2.12us;	slave_if.cable.Current = 	1	;
	#	3us;	slave_if.cable.Current = 	0	;
	#	3.056us;	slave_if.cable.Current = 	1	;
	#	1.104us;	slave_if.cable.Current = 	2	;
	#	1.784us;	slave_if.cable.Current = 	1	;
	#	9.72us;	slave_if.cable.Current = 	2	;
	#	8.112us;	slave_if.cable.Current = 	1	;
	#	6.88us;	slave_if.cable.Current = 	2	;
	#	4.952us;	slave_if.cable.Current = 	1	;
	#	4us;	slave_if.cable.Current = 	2	;
	#	1.952us;	slave_if.cable.Current = 	1	;
	#	9.936us;	slave_if.cable.Current = 	2	;
	#	1.56us;	slave_if.cable.Current = 	1	;
	#	1.056us;	slave_if.cable.Current = 	0	;
	#	2.496us;	slave_if.cable.Current = 	1	;
	#	1.112us;	slave_if.cable.Current = 	2	;
	#	1.672us;	slave_if.cable.Current = 	1	;
	#	6.992us;	slave_if.cable.Current = 	2	;
	#	1.56us;	slave_if.cable.Current = 	1	;
	#	1.056us;	slave_if.cable.Current = 	0	;
	#	5.552us;	slave_if.cable.Current = 	1	;
	#	1.112us;	slave_if.cable.Current = 	2	;
	#	1.616us;	slave_if.cable.Current = 	1	;
	#	8.992us;	slave_if.cable.Current = 	0	;
	#	4.056us;	slave_if.cable.Current = 	1	;
	#	2.944us;	slave_if.cable.Current = 	2	;
	#	1.896us;	slave_if.cable.Current = 	1	;
	#	9.936us;	slave_if.cable.Current = 	2	;
	#	2.008us;	slave_if.cable.Current = 	1	;
	#	6us;	slave_if.cable.Current = 	0	;
	#	3.104us;	slave_if.cable.Current = 	1	;
	#	1.168us;	slave_if.cable.Current = 	2	;
	#	1.616us;	slave_if.cable.Current = 	1	;
	#	6.056us;	slave_if.cable.Current = 	0	;
	#	3.944us;	slave_if.cable.Current = 	1	;
	#	2us;	slave_if.cable.Current = 	0	;
	#	3.16us;	slave_if.cable.Current = 	1	;
	#	1.112us;	slave_if.cable.Current = 	2	;
	#	4.672us;	slave_if.cable.Current = 	1	;
	#	8.944us;	slave_if.cable.Current = 	0	;
	#	3.104us;	slave_if.cable.Current = 	1	;
	#	1.168us;	slave_if.cable.Current = 	2	;
	#	1.672us;	slave_if.cable.Current = 	1	;
	#	3us;	slave_if.cable.Current = 	0	;
	#	3.16us;	slave_if.cable.Current = 	1	;
	#	1.112us;	slave_if.cable.Current = 	2	;
	#	1.672us;	slave_if.cable.Current = 	1	;
	#	3us;	slave_if.cable.Current = 	0	;
	#	3.16us;	slave_if.cable.Current = 	1	;
	#	1.112us;	slave_if.cable.Current = 	2	;
	#	4.232us;	slave_if.cable.Current = 	1	;
	#	1.056us;	slave_if.cable.Current = 	0	;
	#	2.552us;	slave_if.cable.Current = 	1	;
	#	1.272us;	slave_if.cable.Current = 	2	;
	#	1.34399us;	slave_if.cable.Current = 	1	;
	#	3.056us;	slave_if.cable.Current = 	0	;
	#	3.272us;	slave_if.cable.Current = 	1	;
	#	1.216us;	slave_if.cable.Current = 	2	;
	#	1.4us;	slave_if.cable.Current = 	1	;
	#	3.056us;	slave_if.cable.Current = 	0	;
	#	7.272us;	slave_if.cable.Current = 	1	;
	#	1.672us;	slave_if.cable.Current = 	0	;
	#	3.328us;	slave_if.cable.Current = 	1	;
	#	1.216us;	slave_if.cable.Current = 	2	;
	#	4.4us;	slave_if.cable.Current = 	1	;
	#	4.216us;	slave_if.cable.Current = 	2	;
	#	1.728us;	slave_if.cable.Current = 	1	;
	#	2.944us;	slave_if.cable.Current = 	0	;
	#	3.328us;	slave_if.cable.Current = 	1	;
	#	1.224us;	slave_if.cable.Current = 	2	;
	#	1.448us;	slave_if.cable.Current = 	1	;
	#	7.216us;	slave_if.cable.Current = 	2	;
	#	1.728us;	slave_if.cable.Current = 	1	;
	#	2.944us;	slave_if.cable.Current = 	0	;
	#	3.328us;	slave_if.cable.Current = 	1	;
	#	1.272us;	slave_if.cable.Current = 	2	;
	#	4.008us;	slave_if.cable.Current = 	1	;
	#	1.056us;	slave_if.cable.Current = 	0	;
	#	3.608us;	slave_if.cable.Current = 	1	;
	#	4.672us;	slave_if.cable.Current = 	0	;
	#	3.272us;	slave_if.cable.Current = 	1	;
	#	1.224us;	slave_if.cable.Current = 	2	;
	#	7.008us;	slave_if.cable.Current = 	1	;
	#	1.056us;	slave_if.cable.Current = 	0	;
	#	3.544us;	slave_if.cable.Current = 	1	;
	#	1.728us;	slave_if.cable.Current = 	0	;
	#	3.328us;	slave_if.cable.Current = 	1	;
	#	1.224us;	slave_if.cable.Current = 	2	;
	#	4.392us;	slave_if.cable.Current = 	1	;
	#	2.944us;	slave_if.cable.Current = 	0	;
	#	4.328us;	slave_if.cable.Current = 	1	;
	#	1.672us;	slave_if.cable.Current = 	0	;
	#	3.328us;	slave_if.cable.Current = 	1	;
	#	1.224us;	slave_if.cable.Current = 	2	;
	#	1.448us;	slave_if.cable.Current = 	1	;
	#	4.216us;	slave_if.cable.Current = 	2	;
	#	4.672us;	slave_if.cable.Current = 	1	;
	#	3.008us;	slave_if.cable.Current = 	0	;
	#	3.32us;	slave_if.cable.Current = 	1	;
	#	1.224us;	slave_if.cable.Current = 	2	;
	#	7.344us;	slave_if.cable.Current = 	1	;
	#	5.944us;	slave_if.cable.Current = 	0	;
	#	3.32us;	slave_if.cable.Current = 	1	;
	#	1.224us;	slave_if.cable.Current = 	2	;
	#	1.4us;	slave_if.cable.Current = 	1	;
	#	4.272us;	slave_if.cable.Current = 	2	;
	#	1.336us;	slave_if.cable.Current = 	1	;
	#	1.056us;	slave_if.cable.Current = 	0	;
	#	3.552us;	slave_if.cable.Current = 	1	;
	#	1.728us;	slave_if.cable.Current = 	0	;
	#	3.328us;	slave_if.cable.Current = 	1	;
	#	1.16us;	slave_if.cable.Current = 	2	;
	#	4.064us;	slave_if.cable.Current = 	1	;
	#	1.112us;	slave_if.cable.Current = 	0	;
	#	6.552us;	slave_if.cable.Current = 	1	;
	#	1.672us;	slave_if.cable.Current = 	0	;
	#	3.328us;	slave_if.cable.Current = 	1	;
	#	1.216us;	slave_if.cable.Current = 	2	;
	#	1.456us;	slave_if.cable.Current = 	1	;
	#	2.832us;	slave_if.cable.Current = 	0	;
	#	4.608us;	slave_if.cable.Current = 	1	;
	#	4.336us;	slave_if.cable.Current = 	0	;
	#	3.552us;	slave_if.cable.Current = 	1	;
	#	1.44us;	slave_if.cable.Current = 	2	;
	#	0.952us;	slave_if.cable.Current = 	1	;
	#	4.608us;	slave_if.cable.Current = 	2	;
	#	1.392us;	slave_if.cable.Current = 	1	;
	#	4.552us;	slave_if.cable.Current = 	2	;
	#	1.056us;	slave_if.cable.Current = 	1	;
	#	1.168us;	slave_if.cable.Current = 	0	;
	#	2.664us;	slave_if.cable.Current = 	1	;
	#	1.384us;	slave_if.cable.Current = 	2	;
	#	1.008us;	slave_if.cable.Current = 	1	;
	#	6.056us;	slave_if.cable.Current = 	0	;
	#	3.44us;	slave_if.cable.Current = 	1	;
	#	1.392us;	slave_if.cable.Current = 	2	;
	#	0.728us;	slave_if.cable.Current = 	1	;
	#	1.216us;	slave_if.cable.Current = 	0	;
	#	2.664us;	slave_if.cable.Current = 	1	;
	#	1.392us;	slave_if.cable.Current = 	2	;
	#	4.056us;	slave_if.cable.Current = 	1	;
	#	7.552us;	slave_if.cable.Current = 	2	;
	#	1.008us;	slave_if.cable.Current = 	1	;
	#	1.168us;	slave_if.cable.Current = 	0	;
	#	2.656us;	slave_if.cable.Current = 	1	;
	#	1.392us;	slave_if.cable.Current = 	2	;
	#	1.064us;	slave_if.cable.Current = 	1	;
	#	3.056us;	slave_if.cable.Current = 	0	;
	#	3.488us;	slave_if.cable.Current = 	1	;
	#	1.336us;	slave_if.cable.Current = 	2	;
	#	3.728us;	slave_if.cable.Current = 	1	;
	#	1.112us;	slave_if.cable.Current = 	0	;
	#	2.712us;	slave_if.cable.Current = 	1	;
	#	1.392us;	slave_if.cable.Current = 	2	;
	#	3.728us;	slave_if.cable.Current = 	1	;
	#	1.112us;	slave_if.cable.Current = 	0	;
	#	2.712us;	slave_if.cable.Current = 	1	;
	#	1.392us;	slave_if.cable.Current = 	2	;
	#	3.784us;	slave_if.cable.Current = 	1	;
	#	1.056us;	slave_if.cable.Current = 	0	;
	#	2.656us;	slave_if.cable.Current = 	1	;
	#	1.392us;	slave_if.cable.Current = 	2	;
	#	1.064us;	slave_if.cable.Current = 	1	;
	#	3.056us;	slave_if.cable.Current = 	0	;
	#	6.432us;	slave_if.cable.Current = 	1	;
	#	1.392us;	slave_if.cable.Current = 	2	;
	#	0.728us;	slave_if.cable.Current = 	1	;
	#	1.168us;	slave_if.cable.Current = 	0	;
	#	2.72us;	slave_if.cable.Current = 	1	;
	#	1.384us;	slave_if.cable.Current = 	2	;
	#	4.12us;	slave_if.cable.Current = 	1	;
	#	4.44us;	slave_if.cable.Current = 	2	;
	#	4.056us;	slave_if.cable.Current = 	1	;
	#	1.112us;	slave_if.cable.Current = 	0	;
	#	3.832us;	slave_if.cable.Current = 	1	;
	#	2.992us;	slave_if.cable.Current = 	2	;
	#	1.008us;	slave_if.cable.Current = 	1	;
	#	1.112us;	slave_if.cable.Current = 	0	;
	#	2.72us;	slave_if.cable.Current = 	1	;
	#	1.608us;	slave_if.cable.Current = 	2	;
	#	0.064us;	slave_if.cable.Current = 	1	;
	#	1.608us;	slave_if.cable.Current = 	0	;

endtask

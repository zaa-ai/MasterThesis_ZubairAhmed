m_config.configuration_subscriber = new("configuration_subscriber", this);

package otp_wrapper_pkg;

	localparam logic [3:0] c_otp_vrr_dat  = 4'b0100;
	localparam int c_instr_otp_write_ctrl = 160;
	localparam int c_instr_otp_write_conf = 161;
	localparam int c_instr_otp_write = 162;
	localparam int c_instr_otp_write_ecc = 163;
	localparam int c_instr_otp_read = 164;
	localparam int c_instr_otp_read_ecc = 165;
	localparam int c_instr_otpbist_ctrl = 166;
	localparam int c_instr_otpbist_conf = 167;
	localparam int c_instr_otpbist_stat = 168;
	localparam int c_instr_otp_write_pulse_conf = 169;
	localparam int c_instr_sfr_sysmode = 193;
	localparam int c_otp_array_size = 4096;
	localparam int c_otp_wl_adr = 12;
	localparam int c_otp_wl_dat = 12;
	localparam int c_otp_wl_ecc = 0;
	localparam int c_otp_wl_word = 12;
	localparam int c_otp_wl_ctrl = 16;
	localparam int c_otp_cpu_dat = 8;
	localparam logic [31:0] c_otp_prog_key  = 32'b10000100100100010011101110101100;
	localparam int c_otp_wl_mpp = 8;
	localparam int c_otp_wl_mrr = 16;
	localparam int c_otp_wl_mr = 8;
	localparam int c_otp_trp_dat = 7;
	localparam int BL_OTPCTRL = 16;
	localparam int BL_OTP_MON = 2;
	localparam int BIT_EN_AUTO = 0;
	localparam int BIT_EN_OTPCP = 1;
	localparam int BIT_EN_VPP = 2;
	localparam int BIT_OTP_CTRL3 = 3;
	localparam int BIT_EN_OTP = 4;
	localparam int BIT_OTP_CTRL5 = 5;
	localparam int BIT_SEL_OTP = 6;
	localparam int BIT_OTP_CTRL7 = 7;
	localparam int BIT_CTRL_CLK = 8;
	localparam int BIT_CTRL_WE = 9;
	localparam int BIT_OTP_MON_LSB = 10;
	localparam int BIT_OTP_MON_MSB = 11;
	localparam int BIT_AUTOINC = 12;
	localparam int BIT_BYPASS = 13;
	localparam int BIT_OTP_CTRL14 = 14;
	localparam int BIT_OTP_CTRL15 = 15;
	localparam int BL_OTP_CONF = 32;
	localparam int BL_OTP_MPP = 8;
	localparam int BL_OTP_MRR = 16;
	localparam int BL_OTP_MR = 8;
	localparam int BIT_OTP_MPP_LSB = 0;
	localparam int BIT_OTP_MPP_MSB = 7;
	localparam int BIT_OTP_MRR_LSB = 8;
	localparam int BIT_OTP_MRR_MSB = 23;
	localparam int BIT_OTP_MR_LSB = 24;
	localparam int BIT_OTP_MR_MSB = 31;
	localparam int BL_OTP_WRITE_CONFIG = 12;
	localparam int BIT_OTP_WRITE_CONFIG_MSB = 11;
	localparam int BIT_OTP_WRITE_CONFIG_LSB = 0;
	localparam int BL_OTPBISTCTRL = 16;
	localparam int BL_MAX_SOAK = 3;
	localparam int BIT_OTP_PGM = 0;
	localparam int BIT_OTP_READ = 1;
	localparam int BIT_SOAK = 2;
	localparam int BIT_BIST_CTRL3 = 3;
	localparam int BIT_EN_SOAK = 4;
	localparam int BIT_STRESS = 5;
	localparam int BIT_SEL_TRP = 6;
	localparam int BIT_SEL_RD = 7;
	localparam int BIT_SEL_MPP = 8;
	localparam int BIT_SEL_MRR = 9;
	localparam int BIT_SEL_MR = 10;
	localparam int BIT_BIST_CTRL11 = 11;
	localparam int BIT_MAX_SOAK_LSB = 12;
	localparam int BIT_MAX_SOAK_MSB = 14;
	localparam int BIT_BIST_CTRL15 = 15;
	localparam int BL_OTPBISTCONF = 16;
	localparam int BL_TRP = 7;
	localparam int BL_RD_MODE = 2;
	localparam int BL_ECCERR_L = 2;
	localparam int BL_ECCERR_H = 2;
	localparam int BIT_TRP_LSB = 0;
	localparam int BIT_TRP_MSB = 6;
	localparam int BIT_BIST_CONF7 = 7;
	localparam int BIT_RD_MODE_LSB = 8;
	localparam int BIT_RD_MODE_MSB = 9;
	localparam int BIT_BIST_CONF10 = 10;
	localparam int BIT_BIST_CONF11 = 11;
	localparam int BIT_ECCERR_L_LSB = 12;
	localparam int BIT_ECCERR_L_MSB = 13;
	localparam int BIT_ECCERR_H_LSB = 14;
	localparam int BIT_ECCERR_H_MSB = 15;
	localparam int BL_OTPBISTSTAT = 16;
	localparam int BL_PROG_BIT = 6;
	localparam int BL_SOAK_PULSE = 4;
	localparam int BIT_PROG_BIT_LSB = 0;
	localparam int BIT_PROG_BIT_MSB = 5;
	localparam int BIT_BIST_STAT6 = 6;
	localparam int BIT_DONE = 7;
	localparam int BIT_SOAK_PULSE_LSB = 8;
	localparam int BIT_SOAK_PULSE_MSB = 11;
	localparam int BIT_BUSY = 12;
	localparam int BIT_FAIL0 = 13;
	localparam int BIT_FAIL1 = 14;
	localparam int BIT_SOAK_STAT = 15;
	typedef struct packed {
		logic ehv;
		logic oe;
		logic sel;
		logic we;
		logic ck;
		logic [7:0] mr;
		logic [11:0] addr;
	} t_cot_bus;
	typedef struct packed {
		logic [11:0] data;
	} t_dot_bus;
	typedef struct packed {
		logic vppen;
		logic vrren;
		logic [7:0] mpp;
		logic [15:0] mrr;
	} t_ccp_bus;
	typedef struct packed {
		logic clkout;
		logic ppclkout;
	} t_dcp_bus;
endpackage


slave_timing[1][0].info_corner          = 1;
slave_timing[1][0].info_temp__j__       = 125;
slave_timing[1][0].info_i__quite_rec__  = 0.006000000;
slave_timing[1][0].info_dtr__ib__       = -1;
slave_timing[1][0].info_i__offset_rec__ = 0.000000000;
slave_timing[1][0].info_i__max_slave__  = 0.023000000;
slave_timing[1][0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][0].info_r__dsi_bus__    = 5.000;

slave_timing[1][0].t_rxd1[0][1] = 1660ns;
slave_timing[1][0].t_rxd1[1][0] = 1661ns;
slave_timing[1][0].t_rxd1[0][2] = 1253ns;
slave_timing[1][0].t_rxd1[2][0] = 1996ns;
slave_timing[1][0].t_rxd2[0][2] = 1964ns;
slave_timing[1][0].t_rxd2[2][0] = 1240ns;
slave_timing[1][0].t_rxd2[1][2] = 1632ns;
slave_timing[1][0].t_rxd2[2][1] = 1630ns;

slave_timing[1][1].info_corner          = 1;
slave_timing[1][1].info_temp__j__       = 125;
slave_timing[1][1].info_i__quite_rec__  = 0.006000000;
slave_timing[1][1].info_dtr__ib__       = -1;
slave_timing[1][1].info_i__offset_rec__ = 0.000000000;
slave_timing[1][1].info_i__max_slave__  = 0.025000000;
slave_timing[1][1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][1].info_r__dsi_bus__    = 5.000;

slave_timing[1][1].t_rxd1[0][1] = 1597ns;
slave_timing[1][1].t_rxd1[1][0] = 1708ns;
slave_timing[1][1].t_rxd1[0][2] = 1217ns;
slave_timing[1][1].t_rxd1[2][0] = 2027ns;
slave_timing[1][1].t_rxd2[0][2] = 1848ns;
slave_timing[1][1].t_rxd2[2][0] = 1319ns;
slave_timing[1][1].t_rxd2[1][2] = 1464ns;
slave_timing[1][1].t_rxd2[2][1] = 1797ns;

slave_timing[1][2].info_corner          = 1;
slave_timing[1][2].info_temp__j__       = 125;
slave_timing[1][2].info_i__quite_rec__  = 0.006000000;
slave_timing[1][2].info_dtr__ib__       = 1;
slave_timing[1][2].info_i__offset_rec__ = 0.000000000;
slave_timing[1][2].info_i__max_slave__  = 0.023000000;
slave_timing[1][2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][2].info_r__dsi_bus__    = 5.000;

slave_timing[1][2].t_rxd1[0][1] = 1715ns;
slave_timing[1][2].t_rxd1[1][0] = 1600ns;
slave_timing[1][2].t_rxd1[0][2] = 1281ns;
slave_timing[1][2].t_rxd1[2][0] = 1950ns;
slave_timing[1][2].t_rxd2[0][2] = 2090ns;
slave_timing[1][2].t_rxd2[2][0] = 1155ns;
slave_timing[1][2].t_rxd2[1][2] = 1806ns;
slave_timing[1][2].t_rxd2[2][1] = 1484ns;

slave_timing[1][3].info_corner          = 1;
slave_timing[1][3].info_temp__j__       = 125;
slave_timing[1][3].info_i__quite_rec__  = 0.006000000;
slave_timing[1][3].info_dtr__ib__       = 1;
slave_timing[1][3].info_i__offset_rec__ = 0.000000000;
slave_timing[1][3].info_i__max_slave__  = 0.025000000;
slave_timing[1][3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][3].info_r__dsi_bus__    = 5.000;

slave_timing[1][3].t_rxd1[0][1] = 1646ns;
slave_timing[1][3].t_rxd1[1][0] = 1648ns;
slave_timing[1][3].t_rxd1[0][2] = 1242ns;
slave_timing[1][3].t_rxd1[2][0] = 1985ns;
slave_timing[1][3].t_rxd2[0][2] = 1942ns;
slave_timing[1][3].t_rxd2[2][0] = 1249ns;
slave_timing[1][3].t_rxd2[1][2] = 1609ns;
slave_timing[1][3].t_rxd2[2][1] = 1647ns;

slave_timing[1][4].info_corner          = 1;
slave_timing[1][4].info_temp__j__       = 125;
slave_timing[1][4].info_i__quite_rec__  = 0.006000000;
slave_timing[1][4].info_dtr__ib__       = -1;
slave_timing[1][4].info_i__offset_rec__ = 0.000000000;
slave_timing[1][4].info_i__max_slave__  = 0.023000000;
slave_timing[1][4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][4].info_r__dsi_bus__    = 5.000;

slave_timing[1][4].t_rxd1[0][1] = 1853ns;
slave_timing[1][4].t_rxd1[1][0] = 1810ns;
slave_timing[1][4].t_rxd1[0][2] = 1411ns;
slave_timing[1][4].t_rxd1[2][0] = 2139ns;
slave_timing[1][4].t_rxd2[0][2] = 2009ns;
slave_timing[1][4].t_rxd2[2][0] = 1277ns;
slave_timing[1][4].t_rxd2[1][2] = 1659ns;
slave_timing[1][4].t_rxd2[2][1] = 1661ns;

slave_timing[1][5].info_corner          = 1;
slave_timing[1][5].info_temp__j__       = 125;
slave_timing[1][5].info_i__quite_rec__  = 0.006000000;
slave_timing[1][5].info_dtr__ib__       = -1;
slave_timing[1][5].info_i__offset_rec__ = 0.000000000;
slave_timing[1][5].info_i__max_slave__  = 0.025000000;
slave_timing[1][5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][5].info_r__dsi_bus__    = 5.000;

slave_timing[1][5].t_rxd1[0][1] = 1783ns;
slave_timing[1][5].t_rxd1[1][0] = 1856ns;
slave_timing[1][5].t_rxd1[0][2] = 1373ns;
slave_timing[1][5].t_rxd1[2][0] = 2169ns;
slave_timing[1][5].t_rxd2[0][2] = 1897ns;
slave_timing[1][5].t_rxd2[2][0] = 1355ns;
slave_timing[1][5].t_rxd2[1][2] = 1491ns;
slave_timing[1][5].t_rxd2[2][1] = 1821ns;

slave_timing[1][6].info_corner          = 1;
slave_timing[1][6].info_temp__j__       = 125;
slave_timing[1][6].info_i__quite_rec__  = 0.006000000;
slave_timing[1][6].info_dtr__ib__       = 1;
slave_timing[1][6].info_i__offset_rec__ = 0.000000000;
slave_timing[1][6].info_i__max_slave__  = 0.023000000;
slave_timing[1][6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][6].info_r__dsi_bus__    = 5.000;

slave_timing[1][6].t_rxd1[0][1] = 1913ns;
slave_timing[1][6].t_rxd1[1][0] = 1748ns;
slave_timing[1][6].t_rxd1[0][2] = 1439ns;
slave_timing[1][6].t_rxd1[2][0] = 2091ns;
slave_timing[1][6].t_rxd2[0][2] = 2130ns;
slave_timing[1][6].t_rxd2[2][0] = 1191ns;
slave_timing[1][6].t_rxd2[1][2] = 1826ns;
slave_timing[1][6].t_rxd2[2][1] = 1513ns;

slave_timing[1][7].info_corner          = 1;
slave_timing[1][7].info_temp__j__       = 125;
slave_timing[1][7].info_i__quite_rec__  = 0.006000000;
slave_timing[1][7].info_dtr__ib__       = 1;
slave_timing[1][7].info_i__offset_rec__ = 0.000000000;
slave_timing[1][7].info_i__max_slave__  = 0.025000000;
slave_timing[1][7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][7].info_r__dsi_bus__    = 5.000;

slave_timing[1][7].t_rxd1[0][1] = 1838ns;
slave_timing[1][7].t_rxd1[1][0] = 1796ns;
slave_timing[1][7].t_rxd1[0][2] = 1398ns;
slave_timing[1][7].t_rxd1[2][0] = 2121ns;
slave_timing[1][7].t_rxd2[0][2] = 1985ns;
slave_timing[1][7].t_rxd2[2][0] = 1281ns;
slave_timing[1][7].t_rxd2[1][2] = 1633ns;
slave_timing[1][7].t_rxd2[2][1] = 1673ns;

slave_timing[1][8].info_corner          = 1;
slave_timing[1][8].info_temp__j__       = 125;
slave_timing[1][8].info_i__quite_rec__  = 0.003000000;
slave_timing[1][8].info_dtr__ib__       = -1;
slave_timing[1][8].info_i__offset_rec__ = 0.000000000;
slave_timing[1][8].info_i__max_slave__  = 0.023000000;
slave_timing[1][8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][8].info_r__dsi_bus__    = 5.000;

slave_timing[1][8].t_rxd1[0][1] = 1634ns;
slave_timing[1][8].t_rxd1[1][0] = 1656ns;
slave_timing[1][8].t_rxd1[0][2] = 1234ns;
slave_timing[1][8].t_rxd1[2][0] = 1986ns;
slave_timing[1][8].t_rxd2[0][2] = 1944ns;
slave_timing[1][8].t_rxd2[2][0] = 1243ns;
slave_timing[1][8].t_rxd2[1][2] = 1614ns;
slave_timing[1][8].t_rxd2[2][1] = 1618ns;

slave_timing[1][9].info_corner          = 1;
slave_timing[1][9].info_temp__j__       = 125;
slave_timing[1][9].info_i__quite_rec__  = 0.003000000;
slave_timing[1][9].info_dtr__ib__       = -1;
slave_timing[1][9].info_i__offset_rec__ = 0.000000000;
slave_timing[1][9].info_i__max_slave__  = 0.025000000;
slave_timing[1][9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][9].info_r__dsi_bus__    = 5.000;

slave_timing[1][9].t_rxd1[0][1] = 1572ns;
slave_timing[1][9].t_rxd1[1][0] = 1700ns;
slave_timing[1][9].t_rxd1[0][2] = 1202ns;
slave_timing[1][9].t_rxd1[2][0] = 2017ns;
slave_timing[1][9].t_rxd2[0][2] = 1834ns;
slave_timing[1][9].t_rxd2[2][0] = 1322ns;
slave_timing[1][9].t_rxd2[1][2] = 1447ns;
slave_timing[1][9].t_rxd2[2][1] = 1803ns;

slave_timing[1][10].info_corner          = 1;
slave_timing[1][10].info_temp__j__       = 125;
slave_timing[1][10].info_i__quite_rec__  = 0.003000000;
slave_timing[1][10].info_dtr__ib__       = 1;
slave_timing[1][10].info_i__offset_rec__ = 0.000000000;
slave_timing[1][10].info_i__max_slave__  = 0.023000000;
slave_timing[1][10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][10].info_r__dsi_bus__    = 5.000;

slave_timing[1][10].t_rxd1[0][1] = 1676ns;
slave_timing[1][10].t_rxd1[1][0] = 1598ns;
slave_timing[1][10].t_rxd1[0][2] = 1254ns;
slave_timing[1][10].t_rxd1[2][0] = 1942ns;
slave_timing[1][10].t_rxd2[0][2] = 2056ns;
slave_timing[1][10].t_rxd2[2][0] = 1159ns;
slave_timing[1][10].t_rxd2[1][2] = 1775ns;
slave_timing[1][10].t_rxd2[2][1] = 1488ns;

slave_timing[1][11].info_corner          = 1;
slave_timing[1][11].info_temp__j__       = 125;
slave_timing[1][11].info_i__quite_rec__  = 0.003000000;
slave_timing[1][11].info_dtr__ib__       = 1;
slave_timing[1][11].info_i__offset_rec__ = 0.000000000;
slave_timing[1][11].info_i__max_slave__  = 0.025000000;
slave_timing[1][11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][11].info_r__dsi_bus__    = 5.000;

slave_timing[1][11].t_rxd1[0][1] = 1608ns;
slave_timing[1][11].t_rxd1[1][0] = 1645ns;
slave_timing[1][11].t_rxd1[0][2] = 1217ns;
slave_timing[1][11].t_rxd1[2][0] = 1972ns;
slave_timing[1][11].t_rxd2[0][2] = 1918ns;
slave_timing[1][11].t_rxd2[2][0] = 1249ns;
slave_timing[1][11].t_rxd2[1][2] = 1582ns;
slave_timing[1][11].t_rxd2[2][1] = 1631ns;

slave_timing[1][12].info_corner          = 1;
slave_timing[1][12].info_temp__j__       = 125;
slave_timing[1][12].info_i__quite_rec__  = 0.003000000;
slave_timing[1][12].info_dtr__ib__       = -1;
slave_timing[1][12].info_i__offset_rec__ = 0.000000000;
slave_timing[1][12].info_i__max_slave__  = 0.023000000;
slave_timing[1][12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][12].info_r__dsi_bus__    = 5.000;

slave_timing[1][12].t_rxd1[0][1] = 1837ns;
slave_timing[1][12].t_rxd1[1][0] = 1802ns;
slave_timing[1][12].t_rxd1[0][2] = 1401ns;
slave_timing[1][12].t_rxd1[2][0] = 2127ns;
slave_timing[1][12].t_rxd2[0][2] = 1988ns;
slave_timing[1][12].t_rxd2[2][0] = 1279ns;
slave_timing[1][12].t_rxd2[1][2] = 1639ns;
slave_timing[1][12].t_rxd2[2][1] = 1665ns;

slave_timing[1][13].info_corner          = 1;
slave_timing[1][13].info_temp__j__       = 125;
slave_timing[1][13].info_i__quite_rec__  = 0.003000000;
slave_timing[1][13].info_dtr__ib__       = -1;
slave_timing[1][13].info_i__offset_rec__ = 0.000000000;
slave_timing[1][13].info_i__max_slave__  = 0.025000000;
slave_timing[1][13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][13].info_r__dsi_bus__    = 5.000;

slave_timing[1][13].t_rxd1[0][1] = 1770ns;
slave_timing[1][13].t_rxd1[1][0] = 1850ns;
slave_timing[1][13].t_rxd1[0][2] = 1364ns;
slave_timing[1][13].t_rxd1[2][0] = 2158ns;
slave_timing[1][13].t_rxd2[0][2] = 1879ns;
slave_timing[1][13].t_rxd2[2][0] = 1357ns;
slave_timing[1][13].t_rxd2[1][2] = 1475ns;
slave_timing[1][13].t_rxd2[2][1] = 1830ns;

slave_timing[1][14].info_corner          = 1;
slave_timing[1][14].info_temp__j__       = 125;
slave_timing[1][14].info_i__quite_rec__  = 0.003000000;
slave_timing[1][14].info_dtr__ib__       = 1;
slave_timing[1][14].info_i__offset_rec__ = 0.000000000;
slave_timing[1][14].info_i__max_slave__  = 0.023000000;
slave_timing[1][14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][14].info_r__dsi_bus__    = 5.000;

slave_timing[1][14].t_rxd1[0][1] = 1882ns;
slave_timing[1][14].t_rxd1[1][0] = 1746ns;
slave_timing[1][14].t_rxd1[0][2] = 1422ns;
slave_timing[1][14].t_rxd1[2][0] = 2078ns;
slave_timing[1][14].t_rxd2[0][2] = 2095ns;
slave_timing[1][14].t_rxd2[2][0] = 1189ns;
slave_timing[1][14].t_rxd2[1][2] = 1797ns;
slave_timing[1][14].t_rxd2[2][1] = 1520ns;

slave_timing[1][15].info_corner          = 1;
slave_timing[1][15].info_temp__j__       = 125;
slave_timing[1][15].info_i__quite_rec__  = 0.003000000;
slave_timing[1][15].info_dtr__ib__       = 1;
slave_timing[1][15].info_i__offset_rec__ = 0.000000000;
slave_timing[1][15].info_i__max_slave__  = 0.025000000;
slave_timing[1][15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][15].info_r__dsi_bus__    = 5.000;

slave_timing[1][15].t_rxd1[0][1] = 1810ns;
slave_timing[1][15].t_rxd1[1][0] = 1792ns;
slave_timing[1][15].t_rxd1[0][2] = 1367ns;
slave_timing[1][15].t_rxd1[2][0] = 2110ns;
slave_timing[1][15].t_rxd2[0][2] = 1939ns;
slave_timing[1][15].t_rxd2[2][0] = 1280ns;
slave_timing[1][15].t_rxd2[1][2] = 1606ns;
slave_timing[1][15].t_rxd2[2][1] = 1676ns;

slave_timing[1][16].info_corner          = 1;
slave_timing[1][16].info_temp__j__       = 125;
slave_timing[1][16].info_i__quite_rec__  = 0.000000000;
slave_timing[1][16].info_dtr__ib__       = -1;
slave_timing[1][16].info_i__offset_rec__ = 0.000000000;
slave_timing[1][16].info_i__max_slave__  = 0.023000000;
slave_timing[1][16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][16].info_r__dsi_bus__    = 5.000;

slave_timing[1][16].t_rxd1[0][1] = 1620ns;
slave_timing[1][16].t_rxd1[1][0] = 1632ns;
slave_timing[1][16].t_rxd1[0][2] = 1225ns;
slave_timing[1][16].t_rxd1[2][0] = 1962ns;
slave_timing[1][16].t_rxd2[0][2] = 1935ns;
slave_timing[1][16].t_rxd2[2][0] = 1231ns;
slave_timing[1][16].t_rxd2[1][2] = 1616ns;
slave_timing[1][16].t_rxd2[2][1] = 1618ns;

slave_timing[1][17].info_corner          = 1;
slave_timing[1][17].info_temp__j__       = 125;
slave_timing[1][17].info_i__quite_rec__  = 0.000000000;
slave_timing[1][17].info_dtr__ib__       = -1;
slave_timing[1][17].info_i__offset_rec__ = 0.000000000;
slave_timing[1][17].info_i__max_slave__  = 0.025000000;
slave_timing[1][17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][17].info_r__dsi_bus__    = 5.000;

slave_timing[1][17].t_rxd1[0][1] = 1559ns;
slave_timing[1][17].t_rxd1[1][0] = 1677ns;
slave_timing[1][17].t_rxd1[0][2] = 1191ns;
slave_timing[1][17].t_rxd1[2][0] = 1991ns;
slave_timing[1][17].t_rxd2[0][2] = 1822ns;
slave_timing[1][17].t_rxd2[2][0] = 1308ns;
slave_timing[1][17].t_rxd2[1][2] = 1449ns;
slave_timing[1][17].t_rxd2[2][1] = 1781ns;

slave_timing[1][18].info_corner          = 1;
slave_timing[1][18].info_temp__j__       = 125;
slave_timing[1][18].info_i__quite_rec__  = 0.000000000;
slave_timing[1][18].info_dtr__ib__       = 1;
slave_timing[1][18].info_i__offset_rec__ = 0.000000000;
slave_timing[1][18].info_i__max_slave__  = 0.023000000;
slave_timing[1][18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][18].info_r__dsi_bus__    = 5.000;

slave_timing[1][18].t_rxd1[0][1] = 1680ns;
slave_timing[1][18].t_rxd1[1][0] = 1556ns;
slave_timing[1][18].t_rxd1[0][2] = 1251ns;
slave_timing[1][18].t_rxd1[2][0] = 1898ns;
slave_timing[1][18].t_rxd2[0][2] = 2066ns;
slave_timing[1][18].t_rxd2[2][0] = 1124ns;
slave_timing[1][18].t_rxd2[1][2] = 1801ns;
slave_timing[1][18].t_rxd2[2][1] = 1437ns;

slave_timing[1][19].info_corner          = 1;
slave_timing[1][19].info_temp__j__       = 125;
slave_timing[1][19].info_i__quite_rec__  = 0.000000000;
slave_timing[1][19].info_dtr__ib__       = 1;
slave_timing[1][19].info_i__offset_rec__ = 0.000000000;
slave_timing[1][19].info_i__max_slave__  = 0.025000000;
slave_timing[1][19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][19].info_r__dsi_bus__    = 5.000;

slave_timing[1][19].t_rxd1[0][1] = 1610ns;
slave_timing[1][19].t_rxd1[1][0] = 1603ns;
slave_timing[1][19].t_rxd1[0][2] = 1213ns;
slave_timing[1][19].t_rxd1[2][0] = 1931ns;
slave_timing[1][19].t_rxd2[0][2] = 1917ns;
slave_timing[1][19].t_rxd2[2][0] = 1218ns;
slave_timing[1][19].t_rxd2[1][2] = 1601ns;
slave_timing[1][19].t_rxd2[2][1] = 1600ns;

slave_timing[1][20].info_corner          = 1;
slave_timing[1][20].info_temp__j__       = 125;
slave_timing[1][20].info_i__quite_rec__  = 0.000000000;
slave_timing[1][20].info_dtr__ib__       = -1;
slave_timing[1][20].info_i__offset_rec__ = 0.000000000;
slave_timing[1][20].info_i__max_slave__  = 0.023000000;
slave_timing[1][20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][20].info_r__dsi_bus__    = 5.000;

slave_timing[1][20].t_rxd1[0][1] = 1838ns;
slave_timing[1][20].t_rxd1[1][0] = 1778ns;
slave_timing[1][20].t_rxd1[0][2] = 1401ns;
slave_timing[1][20].t_rxd1[2][0] = 2096ns;
slave_timing[1][20].t_rxd2[0][2] = 1972ns;
slave_timing[1][20].t_rxd2[2][0] = 1262ns;
slave_timing[1][20].t_rxd2[1][2] = 1636ns;
slave_timing[1][20].t_rxd2[2][1] = 1645ns;

slave_timing[1][21].info_corner          = 1;
slave_timing[1][21].info_temp__j__       = 125;
slave_timing[1][21].info_i__quite_rec__  = 0.000000000;
slave_timing[1][21].info_dtr__ib__       = -1;
slave_timing[1][21].info_i__offset_rec__ = 0.000000000;
slave_timing[1][21].info_i__max_slave__  = 0.025000000;
slave_timing[1][21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][21].info_r__dsi_bus__    = 5.000;

slave_timing[1][21].t_rxd1[0][1] = 1772ns;
slave_timing[1][21].t_rxd1[1][0] = 1822ns;
slave_timing[1][21].t_rxd1[0][2] = 1349ns;
slave_timing[1][21].t_rxd1[2][0] = 2125ns;
slave_timing[1][21].t_rxd2[0][2] = 1847ns;
slave_timing[1][21].t_rxd2[2][0] = 1339ns;
slave_timing[1][21].t_rxd2[1][2] = 1473ns;
slave_timing[1][21].t_rxd2[2][1] = 1802ns;

slave_timing[1][22].info_corner          = 1;
slave_timing[1][22].info_temp__j__       = 125;
slave_timing[1][22].info_i__quite_rec__  = 0.000000000;
slave_timing[1][22].info_dtr__ib__       = 1;
slave_timing[1][22].info_i__offset_rec__ = 0.000000000;
slave_timing[1][22].info_i__max_slave__  = 0.023000000;
slave_timing[1][22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][22].info_r__dsi_bus__    = 5.000;

slave_timing[1][22].t_rxd1[0][1] = 1911ns;
slave_timing[1][22].t_rxd1[1][0] = 1702ns;
slave_timing[1][22].t_rxd1[0][2] = 1435ns;
slave_timing[1][22].t_rxd1[2][0] = 2032ns;
slave_timing[1][22].t_rxd2[0][2] = 2096ns;
slave_timing[1][22].t_rxd2[2][0] = 1153ns;
slave_timing[1][22].t_rxd2[1][2] = 1819ns;
slave_timing[1][22].t_rxd2[2][1] = 1443ns;

slave_timing[1][23].info_corner          = 1;
slave_timing[1][23].info_temp__j__       = 125;
slave_timing[1][23].info_i__quite_rec__  = 0.000000000;
slave_timing[1][23].info_dtr__ib__       = 1;
slave_timing[1][23].info_i__offset_rec__ = 0.000000000;
slave_timing[1][23].info_i__max_slave__  = 0.025000000;
slave_timing[1][23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][23].info_r__dsi_bus__    = 5.000;

slave_timing[1][23].t_rxd1[0][1] = 1834ns;
slave_timing[1][23].t_rxd1[1][0] = 1747ns;
slave_timing[1][23].t_rxd1[0][2] = 1395ns;
slave_timing[1][23].t_rxd1[2][0] = 2065ns;
slave_timing[1][23].t_rxd2[0][2] = 1952ns;
slave_timing[1][23].t_rxd2[2][0] = 1248ns;
slave_timing[1][23].t_rxd2[1][2] = 1624ns;
slave_timing[1][23].t_rxd2[2][1] = 1623ns;

slave_timing[1][24].info_corner          = 1;
slave_timing[1][24].info_temp__j__       = 125;
slave_timing[1][24].info_i__quite_rec__  = 0.040000000;
slave_timing[1][24].info_dtr__ib__       = -1;
slave_timing[1][24].info_i__offset_rec__ = 0.000000000;
slave_timing[1][24].info_i__max_slave__  = 0.023000000;
slave_timing[1][24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][24].info_r__dsi_bus__    = 5.000;

slave_timing[1][24].t_rxd1[0][1] = 1658ns;
slave_timing[1][24].t_rxd1[1][0] = 1658ns;
slave_timing[1][24].t_rxd1[0][2] = 1240ns;
slave_timing[1][24].t_rxd1[2][0] = 1993ns;
slave_timing[1][24].t_rxd2[0][2] = 1954ns;
slave_timing[1][24].t_rxd2[2][0] = 1244ns;
slave_timing[1][24].t_rxd2[1][2] = 1637ns;
slave_timing[1][24].t_rxd2[2][1] = 1637ns;

slave_timing[1][25].info_corner          = 1;
slave_timing[1][25].info_temp__j__       = 125;
slave_timing[1][25].info_i__quite_rec__  = 0.040000000;
slave_timing[1][25].info_dtr__ib__       = -1;
slave_timing[1][25].info_i__offset_rec__ = 0.000000000;
slave_timing[1][25].info_i__max_slave__  = 0.025000000;
slave_timing[1][25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][25].info_r__dsi_bus__    = 5.000;

slave_timing[1][25].t_rxd1[0][1] = 1594ns;
slave_timing[1][25].t_rxd1[1][0] = 1706ns;
slave_timing[1][25].t_rxd1[0][2] = 1208ns;
slave_timing[1][25].t_rxd1[2][0] = 2041ns;
slave_timing[1][25].t_rxd2[0][2] = 1845ns;
slave_timing[1][25].t_rxd2[2][0] = 1334ns;
slave_timing[1][25].t_rxd2[1][2] = 1467ns;
slave_timing[1][25].t_rxd2[2][1] = 1802ns;

slave_timing[1][26].info_corner          = 1;
slave_timing[1][26].info_temp__j__       = 125;
slave_timing[1][26].info_i__quite_rec__  = 0.040000000;
slave_timing[1][26].info_dtr__ib__       = 1;
slave_timing[1][26].info_i__offset_rec__ = 0.000000000;
slave_timing[1][26].info_i__max_slave__  = 0.023000000;
slave_timing[1][26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][26].info_r__dsi_bus__    = 5.000;

slave_timing[1][26].t_rxd1[0][1] = 1699ns;
slave_timing[1][26].t_rxd1[1][0] = 1615ns;
slave_timing[1][26].t_rxd1[0][2] = 1271ns;
slave_timing[1][26].t_rxd1[2][0] = 1962ns;
slave_timing[1][26].t_rxd2[0][2] = 2082ns;
slave_timing[1][26].t_rxd2[2][0] = 1170ns;
slave_timing[1][26].t_rxd2[1][2] = 1787ns;
slave_timing[1][26].t_rxd2[2][1] = 1498ns;

slave_timing[1][27].info_corner          = 1;
slave_timing[1][27].info_temp__j__       = 125;
slave_timing[1][27].info_i__quite_rec__  = 0.040000000;
slave_timing[1][27].info_dtr__ib__       = 1;
slave_timing[1][27].info_i__offset_rec__ = 0.000000000;
slave_timing[1][27].info_i__max_slave__  = 0.025000000;
slave_timing[1][27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][27].info_r__dsi_bus__    = 5.000;

slave_timing[1][27].t_rxd1[0][1] = 1630ns;
slave_timing[1][27].t_rxd1[1][0] = 1662ns;
slave_timing[1][27].t_rxd1[0][2] = 1235ns;
slave_timing[1][27].t_rxd1[2][0] = 1996ns;
slave_timing[1][27].t_rxd2[0][2] = 1941ns;
slave_timing[1][27].t_rxd2[2][0] = 1260ns;
slave_timing[1][27].t_rxd2[1][2] = 1594ns;
slave_timing[1][27].t_rxd2[2][1] = 1673ns;

slave_timing[1][28].info_corner          = 1;
slave_timing[1][28].info_temp__j__       = 125;
slave_timing[1][28].info_i__quite_rec__  = 0.040000000;
slave_timing[1][28].info_dtr__ib__       = -1;
slave_timing[1][28].info_i__offset_rec__ = 0.000000000;
slave_timing[1][28].info_i__max_slave__  = 0.023000000;
slave_timing[1][28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][28].info_r__dsi_bus__    = 5.000;

slave_timing[1][28].t_rxd1[0][1] = 1743ns;
slave_timing[1][28].t_rxd1[1][0] = 1779ns;
slave_timing[1][28].t_rxd1[0][2] = 1337ns;
slave_timing[1][28].t_rxd1[2][0] = 2100ns;
slave_timing[1][28].t_rxd2[0][2] = 1996ns;
slave_timing[1][28].t_rxd2[2][0] = 1293ns;
slave_timing[1][28].t_rxd2[1][2] = 1656ns;
slave_timing[1][28].t_rxd2[2][1] = 1686ns;

slave_timing[1][29].info_corner          = 1;
slave_timing[1][29].info_temp__j__       = 125;
slave_timing[1][29].info_i__quite_rec__  = 0.040000000;
slave_timing[1][29].info_dtr__ib__       = -1;
slave_timing[1][29].info_i__offset_rec__ = 0.000000000;
slave_timing[1][29].info_i__max_slave__  = 0.025000000;
slave_timing[1][29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][29].info_r__dsi_bus__    = 5.000;

slave_timing[1][29].t_rxd1[0][1] = 1681ns;
slave_timing[1][29].t_rxd1[1][0] = 1822ns;
slave_timing[1][29].t_rxd1[0][2] = 1302ns;
slave_timing[1][29].t_rxd1[2][0] = 2129ns;
slave_timing[1][29].t_rxd2[0][2] = 1891ns;
slave_timing[1][29].t_rxd2[2][0] = 1365ns;
slave_timing[1][29].t_rxd2[1][2] = 1514ns;
slave_timing[1][29].t_rxd2[2][1] = 1821ns;

slave_timing[1][30].info_corner          = 1;
slave_timing[1][30].info_temp__j__       = 125;
slave_timing[1][30].info_i__quite_rec__  = 0.040000000;
slave_timing[1][30].info_dtr__ib__       = 1;
slave_timing[1][30].info_i__offset_rec__ = 0.000000000;
slave_timing[1][30].info_i__max_slave__  = 0.023000000;
slave_timing[1][30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][30].info_r__dsi_bus__    = 5.000;

slave_timing[1][30].t_rxd1[0][1] = 1807ns;
slave_timing[1][30].t_rxd1[1][0] = 1709ns;
slave_timing[1][30].t_rxd1[0][2] = 1369ns;
slave_timing[1][30].t_rxd1[2][0] = 2054ns;
slave_timing[1][30].t_rxd2[0][2] = 2117ns;
slave_timing[1][30].t_rxd2[2][0] = 1212ns;
slave_timing[1][30].t_rxd2[1][2] = 1824ns;
slave_timing[1][30].t_rxd2[2][1] = 1519ns;

slave_timing[1][31].info_corner          = 1;
slave_timing[1][31].info_temp__j__       = 125;
slave_timing[1][31].info_i__quite_rec__  = 0.040000000;
slave_timing[1][31].info_dtr__ib__       = 1;
slave_timing[1][31].info_i__offset_rec__ = 0.000000000;
slave_timing[1][31].info_i__max_slave__  = 0.025000000;
slave_timing[1][31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][31].info_r__dsi_bus__    = 5.000;

slave_timing[1][31].t_rxd1[0][1] = 1737ns;
slave_timing[1][31].t_rxd1[1][0] = 1755ns;
slave_timing[1][31].t_rxd1[0][2] = 1331ns;
slave_timing[1][31].t_rxd1[2][0] = 2084ns;
slave_timing[1][31].t_rxd2[0][2] = 1985ns;
slave_timing[1][31].t_rxd2[2][0] = 1296ns;
slave_timing[1][31].t_rxd2[1][2] = 1636ns;
slave_timing[1][31].t_rxd2[2][1] = 1698ns;

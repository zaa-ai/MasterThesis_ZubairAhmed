/* ###   interface instances   ###################################################### */

TEST_WS_TMR_SEL_WS_if TEST_WS_TMR_SEL_WS (); 
TEST_WS_TMR_VAL_WS_if TEST_WS_TMR_VAL_WS (); 



**------------------------------------------------
** Main
**------------------------------------------------

.subckt top vsup_p hsin0_p hsin1_p hsout0_p hsout1_p
+gnd

.ends

**------------------------------------------------
**------------------------------------------------

/**
 * Interface: sequence_if
 */
interface sequence_if;
	
	int sequence_count = 0;
	string current_sequence;
	
endinterface




slave_timing[0][224+0].info_corner          = 4;
slave_timing[0][224+0].info_temp__j__       = -40;
slave_timing[0][224+0].info_i__quite_rec__  = 0.006000000;
slave_timing[0][224+0].info_dtr__ib__       = -1;
slave_timing[0][224+0].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+0].info_i__max_slave__  = 0.023000000;
slave_timing[0][224+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][224+0].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+0].t_rxd1[0][1] = 1139ns;
slave_timing[0][224+0].t_rxd1[1][0] = 1131ns;
slave_timing[0][224+0].t_rxd1[0][2] = 832ns;
slave_timing[0][224+0].t_rxd1[2][0] = 1435ns;
slave_timing[0][224+0].t_rxd2[0][2] = 1427ns;
slave_timing[0][224+0].t_rxd2[2][0] = 824ns;
slave_timing[0][224+0].t_rxd2[1][2] = 1123ns;
slave_timing[0][224+0].t_rxd2[2][1] = 1112ns;

slave_timing[0][224+1].info_corner          = 4;
slave_timing[0][224+1].info_temp__j__       = -40;
slave_timing[0][224+1].info_i__quite_rec__  = 0.006000000;
slave_timing[0][224+1].info_dtr__ib__       = -1;
slave_timing[0][224+1].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+1].info_i__max_slave__  = 0.025000000;
slave_timing[0][224+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][224+1].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+1].t_rxd1[0][1] = 1086ns;
slave_timing[0][224+1].t_rxd1[1][0] = 1169ns;
slave_timing[0][224+1].t_rxd1[0][2] = 804ns;
slave_timing[0][224+1].t_rxd1[2][0] = 1470ns;
slave_timing[0][224+1].t_rxd2[0][2] = 1315ns;
slave_timing[0][224+1].t_rxd2[2][0] = 881ns;
slave_timing[0][224+1].t_rxd2[1][2] = 987ns;
slave_timing[0][224+1].t_rxd2[2][1] = 1254ns;

slave_timing[0][224+2].info_corner          = 4;
slave_timing[0][224+2].info_temp__j__       = -40;
slave_timing[0][224+2].info_i__quite_rec__  = 0.006000000;
slave_timing[0][224+2].info_dtr__ib__       = 1;
slave_timing[0][224+2].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+2].info_i__max_slave__  = 0.023000000;
slave_timing[0][224+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][224+2].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+2].t_rxd1[0][1] = 1169ns;
slave_timing[0][224+2].t_rxd1[1][0] = 1108ns;
slave_timing[0][224+2].t_rxd1[0][2] = 842ns;
slave_timing[0][224+2].t_rxd1[2][0] = 1415ns;
slave_timing[0][224+2].t_rxd2[0][2] = 1515ns;
slave_timing[0][224+2].t_rxd2[2][0] = 783ns;
slave_timing[0][224+2].t_rxd2[1][2] = 1224ns;
slave_timing[0][224+2].t_rxd2[2][1] = 1032ns;

slave_timing[0][224+3].info_corner          = 4;
slave_timing[0][224+3].info_temp__j__       = -40;
slave_timing[0][224+3].info_i__quite_rec__  = 0.006000000;
slave_timing[0][224+3].info_dtr__ib__       = 1;
slave_timing[0][224+3].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+3].info_i__max_slave__  = 0.025000000;
slave_timing[0][224+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][224+3].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+3].t_rxd1[0][1] = 1112ns;
slave_timing[0][224+3].t_rxd1[1][0] = 1149ns;
slave_timing[0][224+3].t_rxd1[0][2] = 819ns;
slave_timing[0][224+3].t_rxd1[2][0] = 1451ns;
slave_timing[0][224+3].t_rxd2[0][2] = 1381ns;
slave_timing[0][224+3].t_rxd2[2][0] = 848ns;
slave_timing[0][224+3].t_rxd2[1][2] = 1070ns;
slave_timing[0][224+3].t_rxd2[2][1] = 1162ns;

slave_timing[0][224+4].info_corner          = 4;
slave_timing[0][224+4].info_temp__j__       = -40;
slave_timing[0][224+4].info_i__quite_rec__  = 0.006000000;
slave_timing[0][224+4].info_dtr__ib__       = -1;
slave_timing[0][224+4].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+4].info_i__max_slave__  = 0.023000000;
slave_timing[0][224+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][224+4].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+4].t_rxd1[0][1] = 1218ns;
slave_timing[0][224+4].t_rxd1[1][0] = 1202ns;
slave_timing[0][224+4].t_rxd1[0][2] = 887ns;
slave_timing[0][224+4].t_rxd1[2][0] = 1502ns;
slave_timing[0][224+4].t_rxd2[0][2] = 1455ns;
slave_timing[0][224+4].t_rxd2[2][0] = 844ns;
slave_timing[0][224+4].t_rxd2[1][2] = 1134ns;
slave_timing[0][224+4].t_rxd2[2][1] = 1125ns;

slave_timing[0][224+5].info_corner          = 4;
slave_timing[0][224+5].info_temp__j__       = -40;
slave_timing[0][224+5].info_i__quite_rec__  = 0.006000000;
slave_timing[0][224+5].info_dtr__ib__       = -1;
slave_timing[0][224+5].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+5].info_i__max_slave__  = 0.025000000;
slave_timing[0][224+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][224+5].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+5].t_rxd1[0][1] = 1161ns;
slave_timing[0][224+5].t_rxd1[1][0] = 1242ns;
slave_timing[0][224+5].t_rxd1[0][2] = 860ns;
slave_timing[0][224+5].t_rxd1[2][0] = 1534ns;
slave_timing[0][224+5].t_rxd2[0][2] = 1343ns;
slave_timing[0][224+5].t_rxd2[2][0] = 900ns;
slave_timing[0][224+5].t_rxd2[1][2] = 1002ns;
slave_timing[0][224+5].t_rxd2[2][1] = 1262ns;

slave_timing[0][224+6].info_corner          = 4;
slave_timing[0][224+6].info_temp__j__       = -40;
slave_timing[0][224+6].info_i__quite_rec__  = 0.006000000;
slave_timing[0][224+6].info_dtr__ib__       = 1;
slave_timing[0][224+6].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+6].info_i__max_slave__  = 0.023000000;
slave_timing[0][224+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][224+6].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+6].t_rxd1[0][1] = 1242ns;
slave_timing[0][224+6].t_rxd1[1][0] = 1176ns;
slave_timing[0][224+6].t_rxd1[0][2] = 898ns;
slave_timing[0][224+6].t_rxd1[2][0] = 1477ns;
slave_timing[0][224+6].t_rxd2[0][2] = 1544ns;
slave_timing[0][224+6].t_rxd2[2][0] = 801ns;
slave_timing[0][224+6].t_rxd2[1][2] = 1233ns;
slave_timing[0][224+6].t_rxd2[2][1] = 1043ns;

slave_timing[0][224+7].info_corner          = 4;
slave_timing[0][224+7].info_temp__j__       = -40;
slave_timing[0][224+7].info_i__quite_rec__  = 0.006000000;
slave_timing[0][224+7].info_dtr__ib__       = 1;
slave_timing[0][224+7].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+7].info_i__max_slave__  = 0.025000000;
slave_timing[0][224+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][224+7].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+7].t_rxd1[0][1] = 1184ns;
slave_timing[0][224+7].t_rxd1[1][0] = 1216ns;
slave_timing[0][224+7].t_rxd1[0][2] = 868ns;
slave_timing[0][224+7].t_rxd1[2][0] = 1511ns;
slave_timing[0][224+7].t_rxd2[0][2] = 1405ns;
slave_timing[0][224+7].t_rxd2[2][0] = 864ns;
slave_timing[0][224+7].t_rxd2[1][2] = 1082ns;
slave_timing[0][224+7].t_rxd2[2][1] = 1172ns;

slave_timing[0][224+8].info_corner          = 4;
slave_timing[0][224+8].info_temp__j__       = -40;
slave_timing[0][224+8].info_i__quite_rec__  = 0.003000000;
slave_timing[0][224+8].info_dtr__ib__       = -1;
slave_timing[0][224+8].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+8].info_i__max_slave__  = 0.023000000;
slave_timing[0][224+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][224+8].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+8].t_rxd1[0][1] = 1129ns;
slave_timing[0][224+8].t_rxd1[1][0] = 1140ns;
slave_timing[0][224+8].t_rxd1[0][2] = 827ns;
slave_timing[0][224+8].t_rxd1[2][0] = 1449ns;
slave_timing[0][224+8].t_rxd2[0][2] = 1417ns;
slave_timing[0][224+8].t_rxd2[2][0] = 829ns;
slave_timing[0][224+8].t_rxd2[1][2] = 1115ns;
slave_timing[0][224+8].t_rxd2[2][1] = 1118ns;

slave_timing[0][224+9].info_corner          = 4;
slave_timing[0][224+9].info_temp__j__       = -40;
slave_timing[0][224+9].info_i__quite_rec__  = 0.003000000;
slave_timing[0][224+9].info_dtr__ib__       = -1;
slave_timing[0][224+9].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+9].info_i__max_slave__  = 0.025000000;
slave_timing[0][224+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][224+9].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+9].t_rxd1[0][1] = 1079ns;
slave_timing[0][224+9].t_rxd1[1][0] = 1178ns;
slave_timing[0][224+9].t_rxd1[0][2] = 800ns;
slave_timing[0][224+9].t_rxd1[2][0] = 1480ns;
slave_timing[0][224+9].t_rxd2[0][2] = 1307ns;
slave_timing[0][224+9].t_rxd2[2][0] = 884ns;
slave_timing[0][224+9].t_rxd2[1][2] = 981ns;
slave_timing[0][224+9].t_rxd2[2][1] = 1258ns;

slave_timing[0][224+10].info_corner          = 4;
slave_timing[0][224+10].info_temp__j__       = -40;
slave_timing[0][224+10].info_i__quite_rec__  = 0.003000000;
slave_timing[0][224+10].info_dtr__ib__       = 1;
slave_timing[0][224+10].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+10].info_i__max_slave__  = 0.023000000;
slave_timing[0][224+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][224+10].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+10].t_rxd1[0][1] = 1162ns;
slave_timing[0][224+10].t_rxd1[1][0] = 1114ns;
slave_timing[0][224+10].t_rxd1[0][2] = 840ns;
slave_timing[0][224+10].t_rxd1[2][0] = 1420ns;
slave_timing[0][224+10].t_rxd2[0][2] = 1508ns;
slave_timing[0][224+10].t_rxd2[2][0] = 785ns;
slave_timing[0][224+10].t_rxd2[1][2] = 1218ns;
slave_timing[0][224+10].t_rxd2[2][1] = 1033ns;

slave_timing[0][224+11].info_corner          = 4;
slave_timing[0][224+11].info_temp__j__       = -40;
slave_timing[0][224+11].info_i__quite_rec__  = 0.003000000;
slave_timing[0][224+11].info_dtr__ib__       = 1;
slave_timing[0][224+11].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+11].info_i__max_slave__  = 0.025000000;
slave_timing[0][224+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][224+11].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+11].t_rxd1[0][1] = 1105ns;
slave_timing[0][224+11].t_rxd1[1][0] = 1153ns;
slave_timing[0][224+11].t_rxd1[0][2] = 815ns;
slave_timing[0][224+11].t_rxd1[2][0] = 1457ns;
slave_timing[0][224+11].t_rxd2[0][2] = 1374ns;
slave_timing[0][224+11].t_rxd2[2][0] = 850ns;
slave_timing[0][224+11].t_rxd2[1][2] = 1063ns;
slave_timing[0][224+11].t_rxd2[2][1] = 1166ns;

slave_timing[0][224+12].info_corner          = 4;
slave_timing[0][224+12].info_temp__j__       = -40;
slave_timing[0][224+12].info_i__quite_rec__  = 0.003000000;
slave_timing[0][224+12].info_dtr__ib__       = -1;
slave_timing[0][224+12].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+12].info_i__max_slave__  = 0.023000000;
slave_timing[0][224+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][224+12].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+12].t_rxd1[0][1] = 1210ns;
slave_timing[0][224+12].t_rxd1[1][0] = 1215ns;
slave_timing[0][224+12].t_rxd1[0][2] = 883ns;
slave_timing[0][224+12].t_rxd1[2][0] = 1514ns;
slave_timing[0][224+12].t_rxd2[0][2] = 1445ns;
slave_timing[0][224+12].t_rxd2[2][0] = 845ns;
slave_timing[0][224+12].t_rxd2[1][2] = 1125ns;
slave_timing[0][224+12].t_rxd2[2][1] = 1129ns;

slave_timing[0][224+13].info_corner          = 4;
slave_timing[0][224+13].info_temp__j__       = -40;
slave_timing[0][224+13].info_i__quite_rec__  = 0.003000000;
slave_timing[0][224+13].info_dtr__ib__       = -1;
slave_timing[0][224+13].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+13].info_i__max_slave__  = 0.025000000;
slave_timing[0][224+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][224+13].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+13].t_rxd1[0][1] = 1157ns;
slave_timing[0][224+13].t_rxd1[1][0] = 1253ns;
slave_timing[0][224+13].t_rxd1[0][2] = 856ns;
slave_timing[0][224+13].t_rxd1[2][0] = 1546ns;
slave_timing[0][224+13].t_rxd2[0][2] = 1335ns;
slave_timing[0][224+13].t_rxd2[2][0] = 901ns;
slave_timing[0][224+13].t_rxd2[1][2] = 995ns;
slave_timing[0][224+13].t_rxd2[2][1] = 1269ns;

slave_timing[0][224+14].info_corner          = 4;
slave_timing[0][224+14].info_temp__j__       = -40;
slave_timing[0][224+14].info_i__quite_rec__  = 0.003000000;
slave_timing[0][224+14].info_dtr__ib__       = 1;
slave_timing[0][224+14].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+14].info_i__max_slave__  = 0.023000000;
slave_timing[0][224+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][224+14].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+14].t_rxd1[0][1] = 1239ns;
slave_timing[0][224+14].t_rxd1[1][0] = 1183ns;
slave_timing[0][224+14].t_rxd1[0][2] = 893ns;
slave_timing[0][224+14].t_rxd1[2][0] = 1485ns;
slave_timing[0][224+14].t_rxd2[0][2] = 1533ns;
slave_timing[0][224+14].t_rxd2[2][0] = 803ns;
slave_timing[0][224+14].t_rxd2[1][2] = 1222ns;
slave_timing[0][224+14].t_rxd2[2][1] = 1044ns;

slave_timing[0][224+15].info_corner          = 4;
slave_timing[0][224+15].info_temp__j__       = -40;
slave_timing[0][224+15].info_i__quite_rec__  = 0.003000000;
slave_timing[0][224+15].info_dtr__ib__       = 1;
slave_timing[0][224+15].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+15].info_i__max_slave__  = 0.025000000;
slave_timing[0][224+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][224+15].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+15].t_rxd1[0][1] = 1180ns;
slave_timing[0][224+15].t_rxd1[1][0] = 1220ns;
slave_timing[0][224+15].t_rxd1[0][2] = 867ns;
slave_timing[0][224+15].t_rxd1[2][0] = 1516ns;
slave_timing[0][224+15].t_rxd2[0][2] = 1399ns;
slave_timing[0][224+15].t_rxd2[2][0] = 864ns;
slave_timing[0][224+15].t_rxd2[1][2] = 1073ns;
slave_timing[0][224+15].t_rxd2[2][1] = 1174ns;

slave_timing[0][224+16].info_corner          = 4;
slave_timing[0][224+16].info_temp__j__       = -40;
slave_timing[0][224+16].info_i__quite_rec__  = 0.000000000;
slave_timing[0][224+16].info_dtr__ib__       = -1;
slave_timing[0][224+16].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+16].info_i__max_slave__  = 0.023000000;
slave_timing[0][224+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][224+16].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+16].t_rxd1[0][1] = 1143ns;
slave_timing[0][224+16].t_rxd1[1][0] = 1132ns;
slave_timing[0][224+16].t_rxd1[0][2] = 824ns;
slave_timing[0][224+16].t_rxd1[2][0] = 1438ns;
slave_timing[0][224+16].t_rxd2[0][2] = 1412ns;
slave_timing[0][224+16].t_rxd2[2][0] = 825ns;
slave_timing[0][224+16].t_rxd2[1][2] = 1124ns;
slave_timing[0][224+16].t_rxd2[2][1] = 1112ns;

slave_timing[0][224+17].info_corner          = 4;
slave_timing[0][224+17].info_temp__j__       = -40;
slave_timing[0][224+17].info_i__quite_rec__  = 0.000000000;
slave_timing[0][224+17].info_dtr__ib__       = -1;
slave_timing[0][224+17].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+17].info_i__max_slave__  = 0.025000000;
slave_timing[0][224+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][224+17].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+17].t_rxd1[0][1] = 1090ns;
slave_timing[0][224+17].t_rxd1[1][0] = 1168ns;
slave_timing[0][224+17].t_rxd1[0][2] = 800ns;
slave_timing[0][224+17].t_rxd1[2][0] = 1472ns;
slave_timing[0][224+17].t_rxd2[0][2] = 1306ns;
slave_timing[0][224+17].t_rxd2[2][0] = 882ns;
slave_timing[0][224+17].t_rxd2[1][2] = 993ns;
slave_timing[0][224+17].t_rxd2[2][1] = 1254ns;

slave_timing[0][224+18].info_corner          = 4;
slave_timing[0][224+18].info_temp__j__       = -40;
slave_timing[0][224+18].info_i__quite_rec__  = 0.000000000;
slave_timing[0][224+18].info_dtr__ib__       = 1;
slave_timing[0][224+18].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+18].info_i__max_slave__  = 0.023000000;
slave_timing[0][224+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][224+18].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+18].t_rxd1[0][1] = 1154ns;
slave_timing[0][224+18].t_rxd1[1][0] = 1123ns;
slave_timing[0][224+18].t_rxd1[0][2] = 837ns;
slave_timing[0][224+18].t_rxd1[2][0] = 1432ns;
slave_timing[0][224+18].t_rxd2[0][2] = 1501ns;
slave_timing[0][224+18].t_rxd2[2][0] = 790ns;
slave_timing[0][224+18].t_rxd2[1][2] = 1232ns;
slave_timing[0][224+18].t_rxd2[2][1] = 1023ns;

slave_timing[0][224+19].info_corner          = 4;
slave_timing[0][224+19].info_temp__j__       = -40;
slave_timing[0][224+19].info_i__quite_rec__  = 0.000000000;
slave_timing[0][224+19].info_dtr__ib__       = 1;
slave_timing[0][224+19].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+19].info_i__max_slave__  = 0.025000000;
slave_timing[0][224+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][224+19].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+19].t_rxd1[0][1] = 1102ns;
slave_timing[0][224+19].t_rxd1[1][0] = 1161ns;
slave_timing[0][224+19].t_rxd1[0][2] = 812ns;
slave_timing[0][224+19].t_rxd1[2][0] = 1466ns;
slave_timing[0][224+19].t_rxd2[0][2] = 1369ns;
slave_timing[0][224+19].t_rxd2[2][0] = 851ns;
slave_timing[0][224+19].t_rxd2[1][2] = 1057ns;
slave_timing[0][224+19].t_rxd2[2][1] = 1170ns;

slave_timing[0][224+20].info_corner          = 4;
slave_timing[0][224+20].info_temp__j__       = -40;
slave_timing[0][224+20].info_i__quite_rec__  = 0.000000000;
slave_timing[0][224+20].info_dtr__ib__       = -1;
slave_timing[0][224+20].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+20].info_i__max_slave__  = 0.023000000;
slave_timing[0][224+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][224+20].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+20].t_rxd1[0][1] = 1227ns;
slave_timing[0][224+20].t_rxd1[1][0] = 1207ns;
slave_timing[0][224+20].t_rxd1[0][2] = 881ns;
slave_timing[0][224+20].t_rxd1[2][0] = 1506ns;
slave_timing[0][224+20].t_rxd2[0][2] = 1438ns;
slave_timing[0][224+20].t_rxd2[2][0] = 843ns;
slave_timing[0][224+20].t_rxd2[1][2] = 1133ns;
slave_timing[0][224+20].t_rxd2[2][1] = 1122ns;

slave_timing[0][224+21].info_corner          = 4;
slave_timing[0][224+21].info_temp__j__       = -40;
slave_timing[0][224+21].info_i__quite_rec__  = 0.000000000;
slave_timing[0][224+21].info_dtr__ib__       = -1;
slave_timing[0][224+21].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+21].info_i__max_slave__  = 0.025000000;
slave_timing[0][224+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][224+21].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+21].t_rxd1[0][1] = 1149ns;
slave_timing[0][224+21].t_rxd1[1][0] = 1263ns;
slave_timing[0][224+21].t_rxd1[0][2] = 855ns;
slave_timing[0][224+21].t_rxd1[2][0] = 1557ns;
slave_timing[0][224+21].t_rxd2[0][2] = 1332ns;
slave_timing[0][224+21].t_rxd2[2][0] = 909ns;
slave_timing[0][224+21].t_rxd2[1][2] = 989ns;
slave_timing[0][224+21].t_rxd2[2][1] = 1259ns;

slave_timing[0][224+22].info_corner          = 4;
slave_timing[0][224+22].info_temp__j__       = -40;
slave_timing[0][224+22].info_i__quite_rec__  = 0.000000000;
slave_timing[0][224+22].info_dtr__ib__       = 1;
slave_timing[0][224+22].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+22].info_i__max_slave__  = 0.023000000;
slave_timing[0][224+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][224+22].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+22].t_rxd1[0][1] = 1259ns;
slave_timing[0][224+22].t_rxd1[1][0] = 1192ns;
slave_timing[0][224+22].t_rxd1[0][2] = 892ns;
slave_timing[0][224+22].t_rxd1[2][0] = 1495ns;
slave_timing[0][224+22].t_rxd2[0][2] = 1525ns;
slave_timing[0][224+22].t_rxd2[2][0] = 805ns;
slave_timing[0][224+22].t_rxd2[1][2] = 1239ns;
slave_timing[0][224+22].t_rxd2[2][1] = 1032ns;

slave_timing[0][224+23].info_corner          = 4;
slave_timing[0][224+23].info_temp__j__       = -40;
slave_timing[0][224+23].info_i__quite_rec__  = 0.000000000;
slave_timing[0][224+23].info_dtr__ib__       = 1;
slave_timing[0][224+23].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+23].info_i__max_slave__  = 0.025000000;
slave_timing[0][224+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][224+23].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+23].t_rxd1[0][1] = 1178ns;
slave_timing[0][224+23].t_rxd1[1][0] = 1230ns;
slave_timing[0][224+23].t_rxd1[0][2] = 868ns;
slave_timing[0][224+23].t_rxd1[2][0] = 1527ns;
slave_timing[0][224+23].t_rxd2[0][2] = 1395ns;
slave_timing[0][224+23].t_rxd2[2][0] = 865ns;
slave_timing[0][224+23].t_rxd2[1][2] = 1068ns;
slave_timing[0][224+23].t_rxd2[2][1] = 1179ns;

slave_timing[0][224+24].info_corner          = 4;
slave_timing[0][224+24].info_temp__j__       = -40;
slave_timing[0][224+24].info_i__quite_rec__  = 0.040000000;
slave_timing[0][224+24].info_dtr__ib__       = -1;
slave_timing[0][224+24].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+24].info_i__max_slave__  = 0.023000000;
slave_timing[0][224+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][224+24].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+24].t_rxd1[0][1] = 1113ns;
slave_timing[0][224+24].t_rxd1[1][0] = 1136ns;
slave_timing[0][224+24].t_rxd1[0][2] = 820ns;
slave_timing[0][224+24].t_rxd1[2][0] = 1440ns;
slave_timing[0][224+24].t_rxd2[0][2] = 1412ns;
slave_timing[0][224+24].t_rxd2[2][0] = 831ns;
slave_timing[0][224+24].t_rxd2[1][2] = 1112ns;
slave_timing[0][224+24].t_rxd2[2][1] = 1126ns;

slave_timing[0][224+25].info_corner          = 4;
slave_timing[0][224+25].info_temp__j__       = -40;
slave_timing[0][224+25].info_i__quite_rec__  = 0.040000000;
slave_timing[0][224+25].info_dtr__ib__       = -1;
slave_timing[0][224+25].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+25].info_i__max_slave__  = 0.025000000;
slave_timing[0][224+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][224+25].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+25].t_rxd1[0][1] = 1062ns;
slave_timing[0][224+25].t_rxd1[1][0] = 1172ns;
slave_timing[0][224+25].t_rxd1[0][2] = 794ns;
slave_timing[0][224+25].t_rxd1[2][0] = 1473ns;
slave_timing[0][224+25].t_rxd2[0][2] = 1304ns;
slave_timing[0][224+25].t_rxd2[2][0] = 887ns;
slave_timing[0][224+25].t_rxd2[1][2] = 983ns;
slave_timing[0][224+25].t_rxd2[2][1] = 1270ns;

slave_timing[0][224+26].info_corner          = 4;
slave_timing[0][224+26].info_temp__j__       = -40;
slave_timing[0][224+26].info_i__quite_rec__  = 0.040000000;
slave_timing[0][224+26].info_dtr__ib__       = 1;
slave_timing[0][224+26].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+26].info_i__max_slave__  = 0.023000000;
slave_timing[0][224+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][224+26].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+26].t_rxd1[0][1] = 1152ns;
slave_timing[0][224+26].t_rxd1[1][0] = 1104ns;
slave_timing[0][224+26].t_rxd1[0][2] = 836ns;
slave_timing[0][224+26].t_rxd1[2][0] = 1412ns;
slave_timing[0][224+26].t_rxd2[0][2] = 1507ns;
slave_timing[0][224+26].t_rxd2[2][0] = 787ns;
slave_timing[0][224+26].t_rxd2[1][2] = 1219ns;
slave_timing[0][224+26].t_rxd2[2][1] = 1029ns;

slave_timing[0][224+27].info_corner          = 4;
slave_timing[0][224+27].info_temp__j__       = -40;
slave_timing[0][224+27].info_i__quite_rec__  = 0.040000000;
slave_timing[0][224+27].info_dtr__ib__       = 1;
slave_timing[0][224+27].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+27].info_i__max_slave__  = 0.025000000;
slave_timing[0][224+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][224+27].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+27].t_rxd1[0][1] = 1100ns;
slave_timing[0][224+27].t_rxd1[1][0] = 1141ns;
slave_timing[0][224+27].t_rxd1[0][2] = 810ns;
slave_timing[0][224+27].t_rxd1[2][0] = 1446ns;
slave_timing[0][224+27].t_rxd2[0][2] = 1372ns;
slave_timing[0][224+27].t_rxd2[2][0] = 848ns;
slave_timing[0][224+27].t_rxd2[1][2] = 1071ns;
slave_timing[0][224+27].t_rxd2[2][1] = 1164ns;

slave_timing[0][224+28].info_corner          = 4;
slave_timing[0][224+28].info_temp__j__       = -40;
slave_timing[0][224+28].info_i__quite_rec__  = 0.040000000;
slave_timing[0][224+28].info_dtr__ib__       = -1;
slave_timing[0][224+28].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+28].info_i__max_slave__  = 0.023000000;
slave_timing[0][224+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][224+28].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+28].t_rxd1[0][1] = 1150ns;
slave_timing[0][224+28].t_rxd1[1][0] = 1173ns;
slave_timing[0][224+28].t_rxd1[0][2] = 854ns;
slave_timing[0][224+28].t_rxd1[2][0] = 1467ns;
slave_timing[0][224+28].t_rxd2[0][2] = 1425ns;
slave_timing[0][224+28].t_rxd2[2][0] = 849ns;
slave_timing[0][224+28].t_rxd2[1][2] = 1129ns;
slave_timing[0][224+28].t_rxd2[2][1] = 1138ns;

slave_timing[0][224+29].info_corner          = 4;
slave_timing[0][224+29].info_temp__j__       = -40;
slave_timing[0][224+29].info_i__quite_rec__  = 0.040000000;
slave_timing[0][224+29].info_dtr__ib__       = -1;
slave_timing[0][224+29].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+29].info_i__max_slave__  = 0.025000000;
slave_timing[0][224+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][224+29].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+29].t_rxd1[0][1] = 1102ns;
slave_timing[0][224+29].t_rxd1[1][0] = 1206ns;
slave_timing[0][224+29].t_rxd1[0][2] = 830ns;
slave_timing[0][224+29].t_rxd1[2][0] = 1500ns;
slave_timing[0][224+29].t_rxd2[0][2] = 1324ns;
slave_timing[0][224+29].t_rxd2[2][0] = 906ns;
slave_timing[0][224+29].t_rxd2[1][2] = 1003ns;
slave_timing[0][224+29].t_rxd2[2][1] = 1272ns;

slave_timing[0][224+30].info_corner          = 4;
slave_timing[0][224+30].info_temp__j__       = -40;
slave_timing[0][224+30].info_i__quite_rec__  = 0.040000000;
slave_timing[0][224+30].info_dtr__ib__       = 1;
slave_timing[0][224+30].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+30].info_i__max_slave__  = 0.023000000;
slave_timing[0][224+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][224+30].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+30].t_rxd1[0][1] = 1190ns;
slave_timing[0][224+30].t_rxd1[1][0] = 1137ns;
slave_timing[0][224+30].t_rxd1[0][2] = 871ns;
slave_timing[0][224+30].t_rxd1[2][0] = 1436ns;
slave_timing[0][224+30].t_rxd2[0][2] = 1519ns;
slave_timing[0][224+30].t_rxd2[2][0] = 802ns;
slave_timing[0][224+30].t_rxd2[1][2] = 1235ns;
slave_timing[0][224+30].t_rxd2[2][1] = 1047ns;

slave_timing[0][224+31].info_corner          = 4;
slave_timing[0][224+31].info_temp__j__       = -40;
slave_timing[0][224+31].info_i__quite_rec__  = 0.040000000;
slave_timing[0][224+31].info_dtr__ib__       = 1;
slave_timing[0][224+31].info_i__offset_rec__ = 0.000000000;
slave_timing[0][224+31].info_i__max_slave__  = 0.025000000;
slave_timing[0][224+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][224+31].info_r__dsi_bus__    = 5.000;

slave_timing[0][224+31].t_rxd1[0][1] = 1135ns;
slave_timing[0][224+31].t_rxd1[1][0] = 1177ns;
slave_timing[0][224+31].t_rxd1[0][2] = 845ns;
slave_timing[0][224+31].t_rxd1[2][0] = 1468ns;
slave_timing[0][224+31].t_rxd2[0][2] = 1388ns;
slave_timing[0][224+31].t_rxd2[2][0] = 862ns;
slave_timing[0][224+31].t_rxd2[1][2] = 1090ns;
slave_timing[0][224+31].t_rxd2[2][1] = 1171ns;

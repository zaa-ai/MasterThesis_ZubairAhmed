/* ###   interface instances   ###################################################### */

TEST_TOP_TMR_ANA_if TEST_TOP_TMR_ANA (); 
TEST_TOP_TMR_DIG_if TEST_TOP_TMR_DIG (); 
TEST_TOP_TMR_IN_if TEST_TOP_TMR_IN (); 
TEST_TOP_TMR_OUT_CSB_SCK_if TEST_TOP_TMR_OUT_CSB_SCK (); 
TEST_TOP_TMR_OUT_MOSI_MISO_if TEST_TOP_TMR_OUT_MOSI_MISO (); 
TEST_TOP_TMR_OUT_BFWB_SYNCB_if TEST_TOP_TMR_OUT_BFWB_SYNCB (); 
TEST_TOP_TMR_OUT_DAB_INTB_if TEST_TOP_TMR_OUT_DAB_INTB (); 
TEST_TOP_TMR_OUT_RFC_if TEST_TOP_TMR_OUT_RFC (); 



slave_timing[3][96+0].info_corner          = 4;
slave_timing[3][96+0].info_temp__j__       = 125;
slave_timing[3][96+0].info_i__quite_rec__  = 0.006000000;
slave_timing[3][96+0].info_dtr__ib__       = -1;
slave_timing[3][96+0].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+0].info_i__max_slave__  = 0.023000000;
slave_timing[3][96+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][96+0].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+0].t_rxd1[0][1] = 2760ns;
slave_timing[3][96+0].t_rxd1[1][0] = 2698ns;
slave_timing[3][96+0].t_rxd1[0][2] = 2053ns;
slave_timing[3][96+0].t_rxd1[2][0] = 3294ns;
slave_timing[3][96+0].t_rxd2[0][2] = 3359ns;
slave_timing[3][96+0].t_rxd2[2][0] = 2030ns;
slave_timing[3][96+0].t_rxd2[1][2] = 2812ns;
slave_timing[3][96+0].t_rxd2[2][1] = 2684ns;

slave_timing[3][96+1].info_corner          = 4;
slave_timing[3][96+1].info_temp__j__       = 125;
slave_timing[3][96+1].info_i__quite_rec__  = 0.006000000;
slave_timing[3][96+1].info_dtr__ib__       = -1;
slave_timing[3][96+1].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+1].info_i__max_slave__  = 0.025000000;
slave_timing[3][96+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][96+1].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+1].t_rxd1[0][1] = 2648ns;
slave_timing[3][96+1].t_rxd1[1][0] = 2779ns;
slave_timing[3][96+1].t_rxd1[0][2] = 1990ns;
slave_timing[3][96+1].t_rxd1[2][0] = 3348ns;
slave_timing[3][96+1].t_rxd2[0][2] = 3160ns;
slave_timing[3][96+1].t_rxd2[2][0] = 2184ns;
slave_timing[3][96+1].t_rxd2[1][2] = 2515ns;
slave_timing[3][96+1].t_rxd2[2][1] = 2967ns;

slave_timing[3][96+2].info_corner          = 4;
slave_timing[3][96+2].info_temp__j__       = 125;
slave_timing[3][96+2].info_i__quite_rec__  = 0.006000000;
slave_timing[3][96+2].info_dtr__ib__       = 1;
slave_timing[3][96+2].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+2].info_i__max_slave__  = 0.023000000;
slave_timing[3][96+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][96+2].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+2].t_rxd1[0][1] = 2791ns;
slave_timing[3][96+2].t_rxd1[1][0] = 2638ns;
slave_timing[3][96+2].t_rxd1[0][2] = 2062ns;
slave_timing[3][96+2].t_rxd1[2][0] = 3237ns;
slave_timing[3][96+2].t_rxd2[0][2] = 3493ns;
slave_timing[3][96+2].t_rxd2[2][0] = 1909ns;
slave_timing[3][96+2].t_rxd2[1][2] = 3007ns;
slave_timing[3][96+2].t_rxd2[2][1] = 2491ns;

slave_timing[3][96+3].info_corner          = 4;
slave_timing[3][96+3].info_temp__j__       = 125;
slave_timing[3][96+3].info_i__quite_rec__  = 0.006000000;
slave_timing[3][96+3].info_dtr__ib__       = 1;
slave_timing[3][96+3].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+3].info_i__max_slave__  = 0.025000000;
slave_timing[3][96+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][96+3].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+3].t_rxd1[0][1] = 2680ns;
slave_timing[3][96+3].t_rxd1[1][0] = 2715ns;
slave_timing[3][96+3].t_rxd1[0][2] = 1999ns;
slave_timing[3][96+3].t_rxd1[2][0] = 3291ns;
slave_timing[3][96+3].t_rxd2[0][2] = 3260ns;
slave_timing[3][96+3].t_rxd2[2][0] = 2079ns;
slave_timing[3][96+3].t_rxd2[1][2] = 2678ns;
slave_timing[3][96+3].t_rxd2[2][1] = 2777ns;

slave_timing[3][96+4].info_corner          = 4;
slave_timing[3][96+4].info_temp__j__       = 125;
slave_timing[3][96+4].info_i__quite_rec__  = 0.006000000;
slave_timing[3][96+4].info_dtr__ib__       = -1;
slave_timing[3][96+4].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+4].info_i__max_slave__  = 0.023000000;
slave_timing[3][96+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][96+4].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+4].t_rxd1[0][1] = 2931ns;
slave_timing[3][96+4].t_rxd1[1][0] = 2841ns;
slave_timing[3][96+4].t_rxd1[0][2] = 2198ns;
slave_timing[3][96+4].t_rxd1[2][0] = 3423ns;
slave_timing[3][96+4].t_rxd2[0][2] = 3383ns;
slave_timing[3][96+4].t_rxd2[2][0] = 2054ns;
slave_timing[3][96+4].t_rxd2[1][2] = 2835ns;
slave_timing[3][96+4].t_rxd2[2][1] = 2707ns;

slave_timing[3][96+5].info_corner          = 4;
slave_timing[3][96+5].info_temp__j__       = 125;
slave_timing[3][96+5].info_i__quite_rec__  = 0.006000000;
slave_timing[3][96+5].info_dtr__ib__       = -1;
slave_timing[3][96+5].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+5].info_i__max_slave__  = 0.025000000;
slave_timing[3][96+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][96+5].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+5].t_rxd1[0][1] = 2823ns;
slave_timing[3][96+5].t_rxd1[1][0] = 2921ns;
slave_timing[3][96+5].t_rxd1[0][2] = 2147ns;
slave_timing[3][96+5].t_rxd1[2][0] = 3476ns;
slave_timing[3][96+5].t_rxd2[0][2] = 3188ns;
slave_timing[3][96+5].t_rxd2[2][0] = 2206ns;
slave_timing[3][96+5].t_rxd2[1][2] = 2538ns;
slave_timing[3][96+5].t_rxd2[2][1] = 2990ns;

slave_timing[3][96+6].info_corner          = 4;
slave_timing[3][96+6].info_temp__j__       = 125;
slave_timing[3][96+6].info_i__quite_rec__  = 0.006000000;
slave_timing[3][96+6].info_dtr__ib__       = 1;
slave_timing[3][96+6].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+6].info_i__max_slave__  = 0.023000000;
slave_timing[3][96+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][96+6].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+6].t_rxd1[0][1] = 2965ns;
slave_timing[3][96+6].t_rxd1[1][0] = 2766ns;
slave_timing[3][96+6].t_rxd1[0][2] = 2217ns;
slave_timing[3][96+6].t_rxd1[2][0] = 3362ns;
slave_timing[3][96+6].t_rxd2[0][2] = 3514ns;
slave_timing[3][96+6].t_rxd2[2][0] = 1928ns;
slave_timing[3][96+6].t_rxd2[1][2] = 3080ns;
slave_timing[3][96+6].t_rxd2[2][1] = 2478ns;

slave_timing[3][96+7].info_corner          = 4;
slave_timing[3][96+7].info_temp__j__       = 125;
slave_timing[3][96+7].info_i__quite_rec__  = 0.006000000;
slave_timing[3][96+7].info_dtr__ib__       = 1;
slave_timing[3][96+7].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+7].info_i__max_slave__  = 0.025000000;
slave_timing[3][96+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][96+7].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+7].t_rxd1[0][1] = 2841ns;
slave_timing[3][96+7].t_rxd1[1][0] = 2847ns;
slave_timing[3][96+7].t_rxd1[0][2] = 2151ns;
slave_timing[3][96+7].t_rxd1[2][0] = 3416ns;
slave_timing[3][96+7].t_rxd2[0][2] = 3283ns;
slave_timing[3][96+7].t_rxd2[2][0] = 2100ns;
slave_timing[3][96+7].t_rxd2[1][2] = 2739ns;
slave_timing[3][96+7].t_rxd2[2][1] = 2758ns;

slave_timing[3][96+8].info_corner          = 4;
slave_timing[3][96+8].info_temp__j__       = 125;
slave_timing[3][96+8].info_i__quite_rec__  = 0.003000000;
slave_timing[3][96+8].info_dtr__ib__       = -1;
slave_timing[3][96+8].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+8].info_i__max_slave__  = 0.023000000;
slave_timing[3][96+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][96+8].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+8].t_rxd1[0][1] = 2721ns;
slave_timing[3][96+8].t_rxd1[1][0] = 2664ns;
slave_timing[3][96+8].t_rxd1[0][2] = 2024ns;
slave_timing[3][96+8].t_rxd1[2][0] = 3252ns;
slave_timing[3][96+8].t_rxd2[0][2] = 3329ns;
slave_timing[3][96+8].t_rxd2[2][0] = 1998ns;
slave_timing[3][96+8].t_rxd2[1][2] = 2836ns;
slave_timing[3][96+8].t_rxd2[2][1] = 2606ns;

slave_timing[3][96+9].info_corner          = 4;
slave_timing[3][96+9].info_temp__j__       = 125;
slave_timing[3][96+9].info_i__quite_rec__  = 0.003000000;
slave_timing[3][96+9].info_dtr__ib__       = -1;
slave_timing[3][96+9].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+9].info_i__max_slave__  = 0.025000000;
slave_timing[3][96+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][96+9].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+9].t_rxd1[0][1] = 2615ns;
slave_timing[3][96+9].t_rxd1[1][0] = 2747ns;
slave_timing[3][96+9].t_rxd1[0][2] = 1956ns;
slave_timing[3][96+9].t_rxd1[2][0] = 3306ns;
slave_timing[3][96+9].t_rxd2[0][2] = 3129ns;
slave_timing[3][96+9].t_rxd2[2][0] = 2152ns;
slave_timing[3][96+9].t_rxd2[1][2] = 2496ns;
slave_timing[3][96+9].t_rxd2[2][1] = 2919ns;

slave_timing[3][96+10].info_corner          = 4;
slave_timing[3][96+10].info_temp__j__       = 125;
slave_timing[3][96+10].info_i__quite_rec__  = 0.003000000;
slave_timing[3][96+10].info_dtr__ib__       = 1;
slave_timing[3][96+10].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+10].info_i__max_slave__  = 0.023000000;
slave_timing[3][96+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][96+10].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+10].t_rxd1[0][1] = 2777ns;
slave_timing[3][96+10].t_rxd1[1][0] = 2608ns;
slave_timing[3][96+10].t_rxd1[0][2] = 2045ns;
slave_timing[3][96+10].t_rxd1[2][0] = 3202ns;
slave_timing[3][96+10].t_rxd2[0][2] = 3464ns;
slave_timing[3][96+10].t_rxd2[2][0] = 1857ns;
slave_timing[3][96+10].t_rxd2[1][2] = 2996ns;
slave_timing[3][96+10].t_rxd2[2][1] = 2434ns;

slave_timing[3][96+11].info_corner          = 4;
slave_timing[3][96+11].info_temp__j__       = 125;
slave_timing[3][96+11].info_i__quite_rec__  = 0.003000000;
slave_timing[3][96+11].info_dtr__ib__       = 1;
slave_timing[3][96+11].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+11].info_i__max_slave__  = 0.025000000;
slave_timing[3][96+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][96+11].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+11].t_rxd1[0][1] = 2658ns;
slave_timing[3][96+11].t_rxd1[1][0] = 2687ns;
slave_timing[3][96+11].t_rxd1[0][2] = 1978ns;
slave_timing[3][96+11].t_rxd1[2][0] = 3255ns;
slave_timing[3][96+11].t_rxd2[0][2] = 3230ns;
slave_timing[3][96+11].t_rxd2[2][0] = 2031ns;
slave_timing[3][96+11].t_rxd2[1][2] = 2665ns;
slave_timing[3][96+11].t_rxd2[2][1] = 2710ns;

slave_timing[3][96+12].info_corner          = 4;
slave_timing[3][96+12].info_temp__j__       = 125;
slave_timing[3][96+12].info_i__quite_rec__  = 0.003000000;
slave_timing[3][96+12].info_dtr__ib__       = -1;
slave_timing[3][96+12].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+12].info_i__max_slave__  = 0.023000000;
slave_timing[3][96+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][96+12].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+12].t_rxd1[0][1] = 2911ns;
slave_timing[3][96+12].t_rxd1[1][0] = 2810ns;
slave_timing[3][96+12].t_rxd1[0][2] = 2196ns;
slave_timing[3][96+12].t_rxd1[2][0] = 3387ns;
slave_timing[3][96+12].t_rxd2[0][2] = 3351ns;
slave_timing[3][96+12].t_rxd2[2][0] = 2025ns;
slave_timing[3][96+12].t_rxd2[1][2] = 2856ns;
slave_timing[3][96+12].t_rxd2[2][1] = 2626ns;

slave_timing[3][96+13].info_corner          = 4;
slave_timing[3][96+13].info_temp__j__       = 125;
slave_timing[3][96+13].info_i__quite_rec__  = 0.003000000;
slave_timing[3][96+13].info_dtr__ib__       = -1;
slave_timing[3][96+13].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+13].info_i__max_slave__  = 0.025000000;
slave_timing[3][96+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][96+13].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+13].t_rxd1[0][1] = 2802ns;
slave_timing[3][96+13].t_rxd1[1][0] = 2894ns;
slave_timing[3][96+13].t_rxd1[0][2] = 2126ns;
slave_timing[3][96+13].t_rxd1[2][0] = 3436ns;
slave_timing[3][96+13].t_rxd2[0][2] = 3147ns;
slave_timing[3][96+13].t_rxd2[2][0] = 2174ns;
slave_timing[3][96+13].t_rxd2[1][2] = 2523ns;
slave_timing[3][96+13].t_rxd2[2][1] = 2933ns;

slave_timing[3][96+14].info_corner          = 4;
slave_timing[3][96+14].info_temp__j__       = 125;
slave_timing[3][96+14].info_i__quite_rec__  = 0.003000000;
slave_timing[3][96+14].info_dtr__ib__       = 1;
slave_timing[3][96+14].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+14].info_i__max_slave__  = 0.023000000;
slave_timing[3][96+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][96+14].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+14].t_rxd1[0][1] = 2960ns;
slave_timing[3][96+14].t_rxd1[1][0] = 2747ns;
slave_timing[3][96+14].t_rxd1[0][2] = 2210ns;
slave_timing[3][96+14].t_rxd1[2][0] = 3330ns;
slave_timing[3][96+14].t_rxd2[0][2] = 3479ns;
slave_timing[3][96+14].t_rxd2[2][0] = 1877ns;
slave_timing[3][96+14].t_rxd2[1][2] = 3015ns;
slave_timing[3][96+14].t_rxd2[2][1] = 2448ns;

slave_timing[3][96+15].info_corner          = 4;
slave_timing[3][96+15].info_temp__j__       = 125;
slave_timing[3][96+15].info_i__quite_rec__  = 0.003000000;
slave_timing[3][96+15].info_dtr__ib__       = 1;
slave_timing[3][96+15].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+15].info_i__max_slave__  = 0.025000000;
slave_timing[3][96+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][96+15].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+15].t_rxd1[0][1] = 2837ns;
slave_timing[3][96+15].t_rxd1[1][0] = 2826ns;
slave_timing[3][96+15].t_rxd1[0][2] = 2146ns;
slave_timing[3][96+15].t_rxd1[2][0] = 3379ns;
slave_timing[3][96+15].t_rxd2[0][2] = 3248ns;
slave_timing[3][96+15].t_rxd2[2][0] = 2049ns;
slave_timing[3][96+15].t_rxd2[1][2] = 2682ns;
slave_timing[3][96+15].t_rxd2[2][1] = 2728ns;

slave_timing[3][96+16].info_corner          = 4;
slave_timing[3][96+16].info_temp__j__       = 125;
slave_timing[3][96+16].info_i__quite_rec__  = 0.000000000;
slave_timing[3][96+16].info_dtr__ib__       = -1;
slave_timing[3][96+16].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+16].info_i__max_slave__  = 0.023000000;
slave_timing[3][96+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][96+16].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+16].t_rxd1[0][1] = 2700ns;
slave_timing[3][96+16].t_rxd1[1][0] = 2641ns;
slave_timing[3][96+16].t_rxd1[0][2] = 1984ns;
slave_timing[3][96+16].t_rxd1[2][0] = 3215ns;
slave_timing[3][96+16].t_rxd2[0][2] = 3286ns;
slave_timing[3][96+16].t_rxd2[2][0] = 1953ns;
slave_timing[3][96+16].t_rxd2[1][2] = 2765ns;
slave_timing[3][96+16].t_rxd2[2][1] = 2587ns;

slave_timing[3][96+17].info_corner          = 4;
slave_timing[3][96+17].info_temp__j__       = 125;
slave_timing[3][96+17].info_i__quite_rec__  = 0.000000000;
slave_timing[3][96+17].info_dtr__ib__       = -1;
slave_timing[3][96+17].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+17].info_i__max_slave__  = 0.025000000;
slave_timing[3][96+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][96+17].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+17].t_rxd1[0][1] = 2597ns;
slave_timing[3][96+17].t_rxd1[1][0] = 2719ns;
slave_timing[3][96+17].t_rxd1[0][2] = 1943ns;
slave_timing[3][96+17].t_rxd1[2][0] = 3269ns;
slave_timing[3][96+17].t_rxd2[0][2] = 3084ns;
slave_timing[3][96+17].t_rxd2[2][0] = 2107ns;
slave_timing[3][96+17].t_rxd2[1][2] = 2473ns;
slave_timing[3][96+17].t_rxd2[2][1] = 2864ns;

slave_timing[3][96+18].info_corner          = 4;
slave_timing[3][96+18].info_temp__j__       = 125;
slave_timing[3][96+18].info_i__quite_rec__  = 0.000000000;
slave_timing[3][96+18].info_dtr__ib__       = 1;
slave_timing[3][96+18].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+18].info_i__max_slave__  = 0.023000000;
slave_timing[3][96+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][96+18].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+18].t_rxd1[0][1] = 2738ns;
slave_timing[3][96+18].t_rxd1[1][0] = 2576ns;
slave_timing[3][96+18].t_rxd1[0][2] = 2023ns;
slave_timing[3][96+18].t_rxd1[2][0] = 3167ns;
slave_timing[3][96+18].t_rxd2[0][2] = 3425ns;
slave_timing[3][96+18].t_rxd2[2][0] = 1820ns;
slave_timing[3][96+18].t_rxd2[1][2] = 2966ns;
slave_timing[3][96+18].t_rxd2[2][1] = 2383ns;

slave_timing[3][96+19].info_corner          = 4;
slave_timing[3][96+19].info_temp__j__       = 125;
slave_timing[3][96+19].info_i__quite_rec__  = 0.000000000;
slave_timing[3][96+19].info_dtr__ib__       = 1;
slave_timing[3][96+19].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+19].info_i__max_slave__  = 0.025000000;
slave_timing[3][96+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][96+19].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+19].t_rxd1[0][1] = 2629ns;
slave_timing[3][96+19].t_rxd1[1][0] = 2657ns;
slave_timing[3][96+19].t_rxd1[0][2] = 1959ns;
slave_timing[3][96+19].t_rxd1[2][0] = 3222ns;
slave_timing[3][96+19].t_rxd2[0][2] = 3191ns;
slave_timing[3][96+19].t_rxd2[2][0] = 1996ns;
slave_timing[3][96+19].t_rxd2[1][2] = 2636ns;
slave_timing[3][96+19].t_rxd2[2][1] = 2663ns;

slave_timing[3][96+20].info_corner          = 4;
slave_timing[3][96+20].info_temp__j__       = 125;
slave_timing[3][96+20].info_i__quite_rec__  = 0.000000000;
slave_timing[3][96+20].info_dtr__ib__       = -1;
slave_timing[3][96+20].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+20].info_i__max_slave__  = 0.023000000;
slave_timing[3][96+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][96+20].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+20].t_rxd1[0][1] = 2907ns;
slave_timing[3][96+20].t_rxd1[1][0] = 2787ns;
slave_timing[3][96+20].t_rxd1[0][2] = 2193ns;
slave_timing[3][96+20].t_rxd1[2][0] = 3350ns;
slave_timing[3][96+20].t_rxd2[0][2] = 3300ns;
slave_timing[3][96+20].t_rxd2[2][0] = 1976ns;
slave_timing[3][96+20].t_rxd2[1][2] = 2818ns;
slave_timing[3][96+20].t_rxd2[2][1] = 2576ns;

slave_timing[3][96+21].info_corner          = 4;
slave_timing[3][96+21].info_temp__j__       = 125;
slave_timing[3][96+21].info_i__quite_rec__  = 0.000000000;
slave_timing[3][96+21].info_dtr__ib__       = -1;
slave_timing[3][96+21].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+21].info_i__max_slave__  = 0.025000000;
slave_timing[3][96+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][96+21].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+21].t_rxd1[0][1] = 2797ns;
slave_timing[3][96+21].t_rxd1[1][0] = 2860ns;
slave_timing[3][96+21].t_rxd1[0][2] = 2127ns;
slave_timing[3][96+21].t_rxd1[2][0] = 3398ns;
slave_timing[3][96+21].t_rxd2[0][2] = 3102ns;
slave_timing[3][96+21].t_rxd2[2][0] = 2132ns;
slave_timing[3][96+21].t_rxd2[1][2] = 2509ns;
slave_timing[3][96+21].t_rxd2[2][1] = 2844ns;

slave_timing[3][96+22].info_corner          = 4;
slave_timing[3][96+22].info_temp__j__       = 125;
slave_timing[3][96+22].info_i__quite_rec__  = 0.000000000;
slave_timing[3][96+22].info_dtr__ib__       = 1;
slave_timing[3][96+22].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+22].info_i__max_slave__  = 0.023000000;
slave_timing[3][96+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][96+22].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+22].t_rxd1[0][1] = 2945ns;
slave_timing[3][96+22].t_rxd1[1][0] = 2714ns;
slave_timing[3][96+22].t_rxd1[0][2] = 2200ns;
slave_timing[3][96+22].t_rxd1[2][0] = 3298ns;
slave_timing[3][96+22].t_rxd2[0][2] = 3437ns;
slave_timing[3][96+22].t_rxd2[2][0] = 1839ns;
slave_timing[3][96+22].t_rxd2[1][2] = 3034ns;
slave_timing[3][96+22].t_rxd2[2][1] = 2370ns;

slave_timing[3][96+23].info_corner          = 4;
slave_timing[3][96+23].info_temp__j__       = 125;
slave_timing[3][96+23].info_i__quite_rec__  = 0.000000000;
slave_timing[3][96+23].info_dtr__ib__       = 1;
slave_timing[3][96+23].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+23].info_i__max_slave__  = 0.025000000;
slave_timing[3][96+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][96+23].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+23].t_rxd1[0][1] = 2829ns;
slave_timing[3][96+23].t_rxd1[1][0] = 2795ns;
slave_timing[3][96+23].t_rxd1[0][2] = 2136ns;
slave_timing[3][96+23].t_rxd1[2][0] = 3351ns;
slave_timing[3][96+23].t_rxd2[0][2] = 3203ns;
slave_timing[3][96+23].t_rxd2[2][0] = 2016ns;
slave_timing[3][96+23].t_rxd2[1][2] = 2692ns;
slave_timing[3][96+23].t_rxd2[2][1] = 2648ns;

slave_timing[3][96+24].info_corner          = 4;
slave_timing[3][96+24].info_temp__j__       = 125;
slave_timing[3][96+24].info_i__quite_rec__  = 0.040000000;
slave_timing[3][96+24].info_dtr__ib__       = -1;
slave_timing[3][96+24].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+24].info_i__max_slave__  = 0.023000000;
slave_timing[3][96+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][96+24].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+24].t_rxd1[0][1] = 2801ns;
slave_timing[3][96+24].t_rxd1[1][0] = 2747ns;
slave_timing[3][96+24].t_rxd1[0][2] = 2114ns;
slave_timing[3][96+24].t_rxd1[2][0] = 3393ns;
slave_timing[3][96+24].t_rxd2[0][2] = 3634ns;
slave_timing[3][96+24].t_rxd2[2][0] = 2265ns;
slave_timing[3][96+24].t_rxd2[1][2] = 3055ns;
slave_timing[3][96+24].t_rxd2[2][1] = 2967ns;

slave_timing[3][96+25].info_corner          = 4;
slave_timing[3][96+25].info_temp__j__       = 125;
slave_timing[3][96+25].info_i__quite_rec__  = 0.040000000;
slave_timing[3][96+25].info_dtr__ib__       = -1;
slave_timing[3][96+25].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+25].info_i__max_slave__  = 0.025000000;
slave_timing[3][96+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][96+25].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+25].t_rxd1[0][1] = 2700ns;
slave_timing[3][96+25].t_rxd1[1][0] = 2835ns;
slave_timing[3][96+25].t_rxd1[0][2] = 2053ns;
slave_timing[3][96+25].t_rxd1[2][0] = 3451ns;
slave_timing[3][96+25].t_rxd2[0][2] = 3431ns;
slave_timing[3][96+25].t_rxd2[2][0] = 2414ns;
slave_timing[3][96+25].t_rxd2[1][2] = 2748ns;
slave_timing[3][96+25].t_rxd2[2][1] = 3218ns;

slave_timing[3][96+26].info_corner          = 4;
slave_timing[3][96+26].info_temp__j__       = 125;
slave_timing[3][96+26].info_i__quite_rec__  = 0.040000000;
slave_timing[3][96+26].info_dtr__ib__       = 1;
slave_timing[3][96+26].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+26].info_i__max_slave__  = 0.023000000;
slave_timing[3][96+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][96+26].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+26].t_rxd1[0][1] = 2895ns;
slave_timing[3][96+26].t_rxd1[1][0] = 2673ns;
slave_timing[3][96+26].t_rxd1[0][2] = 2164ns;
slave_timing[3][96+26].t_rxd1[2][0] = 3345ns;
slave_timing[3][96+26].t_rxd2[0][2] = 3804ns;
slave_timing[3][96+26].t_rxd2[2][0] = 2136ns;
slave_timing[3][96+26].t_rxd2[1][2] = 3299ns;
slave_timing[3][96+26].t_rxd2[2][1] = 2750ns;

slave_timing[3][96+27].info_corner          = 4;
slave_timing[3][96+27].info_temp__j__       = 125;
slave_timing[3][96+27].info_i__quite_rec__  = 0.040000000;
slave_timing[3][96+27].info_dtr__ib__       = 1;
slave_timing[3][96+27].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+27].info_i__max_slave__  = 0.025000000;
slave_timing[3][96+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][96+27].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+27].t_rxd1[0][1] = 2775ns;
slave_timing[3][96+27].t_rxd1[1][0] = 2768ns;
slave_timing[3][96+27].t_rxd1[0][2] = 2101ns;
slave_timing[3][96+27].t_rxd1[2][0] = 3404ns;
slave_timing[3][96+27].t_rxd2[0][2] = 3561ns;
slave_timing[3][96+27].t_rxd2[2][0] = 2306ns;
slave_timing[3][96+27].t_rxd2[1][2] = 2956ns;
slave_timing[3][96+27].t_rxd2[2][1] = 3045ns;

slave_timing[3][96+28].info_corner          = 4;
slave_timing[3][96+28].info_temp__j__       = 125;
slave_timing[3][96+28].info_i__quite_rec__  = 0.040000000;
slave_timing[3][96+28].info_dtr__ib__       = -1;
slave_timing[3][96+28].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+28].info_i__max_slave__  = 0.023000000;
slave_timing[3][96+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][96+28].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+28].t_rxd1[0][1] = 2875ns;
slave_timing[3][96+28].t_rxd1[1][0] = 3127ns;
slave_timing[3][96+28].t_rxd1[0][2] = 2201ns;
slave_timing[3][96+28].t_rxd1[2][0] = 4164ns;
slave_timing[3][96+28].t_rxd2[0][2] = 4570ns;
slave_timing[3][96+28].t_rxd2[2][0] = 2884ns;
slave_timing[3][96+28].t_rxd2[1][2] = 3910ns;
slave_timing[3][96+28].t_rxd2[2][1] = 3817ns;

slave_timing[3][96+29].info_corner          = 4;
slave_timing[3][96+29].info_temp__j__       = 125;
slave_timing[3][96+29].info_i__quite_rec__  = 0.040000000;
slave_timing[3][96+29].info_dtr__ib__       = -1;
slave_timing[3][96+29].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+29].info_i__max_slave__  = 0.025000000;
slave_timing[3][96+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][96+29].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+29].t_rxd1[0][1] = 2778ns;
slave_timing[3][96+29].t_rxd1[1][0] = 3267ns;
slave_timing[3][96+29].t_rxd1[0][2] = 2144ns;
slave_timing[3][96+29].t_rxd1[2][0] = 4267ns;
slave_timing[3][96+29].t_rxd2[0][2] = 4262ns;
slave_timing[3][96+29].t_rxd2[2][0] = 3079ns;
slave_timing[3][96+29].t_rxd2[1][2] = 3488ns;
slave_timing[3][96+29].t_rxd2[2][1] = 4252ns;

slave_timing[3][96+30].info_corner          = 4;
slave_timing[3][96+30].info_temp__j__       = 125;
slave_timing[3][96+30].info_i__quite_rec__  = 0.040000000;
slave_timing[3][96+30].info_dtr__ib__       = 1;
slave_timing[3][96+30].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+30].info_i__max_slave__  = 0.023000000;
slave_timing[3][96+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][96+30].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+30].t_rxd1[0][1] = 2962ns;
slave_timing[3][96+30].t_rxd1[1][0] = 2968ns;
slave_timing[3][96+30].t_rxd1[0][2] = 2251ns;
slave_timing[3][96+30].t_rxd1[2][0] = 4037ns;
slave_timing[3][96+30].t_rxd2[0][2] = 4835ns;
slave_timing[3][96+30].t_rxd2[2][0] = 2714ns;
slave_timing[3][96+30].t_rxd2[1][2] = 4247ns;
slave_timing[3][96+30].t_rxd2[2][1] = 3507ns;

slave_timing[3][96+31].info_corner          = 4;
slave_timing[3][96+31].info_temp__j__       = 125;
slave_timing[3][96+31].info_i__quite_rec__  = 0.040000000;
slave_timing[3][96+31].info_dtr__ib__       = 1;
slave_timing[3][96+31].info_i__offset_rec__ = 0.000000000;
slave_timing[3][96+31].info_i__max_slave__  = 0.025000000;
slave_timing[3][96+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][96+31].info_r__dsi_bus__    = 5.000;

slave_timing[3][96+31].t_rxd1[0][1] = 2847ns;
slave_timing[3][96+31].t_rxd1[1][0] = 3113ns;
slave_timing[3][96+31].t_rxd1[0][2] = 2188ns;
slave_timing[3][96+31].t_rxd1[2][0] = 4141ns;
slave_timing[3][96+31].t_rxd2[0][2] = 4448ns;
slave_timing[3][96+31].t_rxd2[2][0] = 2931ns;
slave_timing[3][96+31].t_rxd2[1][2] = 3762ns;
slave_timing[3][96+31].t_rxd2[2][1] = 3919ns;

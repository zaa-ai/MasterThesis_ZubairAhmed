/**
 * Package: unit_test_pkg
 * 
 * package for unit testing
 */
package unit_test_pkg;
	import uvm_pkg::*;
	import common_env_pkg::*;
	import project_pkg::*;
	import elip_bus_pkg::*;
	import ECC_pkg::*;
	
	`include "agent_factory.svh"
	`include "top_config.svh"
	`include "top_env.svh"
	`include "top_test.svh"

endpackage



//-----------------------------------------------------------------------------
// Copyright (c) 2023 Elmos SE
// Author     : Eugene - Easy UVM Generator
//
// Description: This file has been generated automatically by Eugene
//				This file should not be modified manually. 
//-----------------------------------------------------------------------------
`ifndef DIGITAL_SIGNAL_MONITOR_SV
`define DIGITAL_SIGNAL_MONITOR_SV

class digital_signal_monitor extends uvm_monitor;

	`uvm_component_utils(digital_signal_monitor)
	
	virtual	digital_signal_if vif;

  	digital_signal_config m_config;

  	uvm_analysis_port #(digital_signal_tr) analysis_port;

  	digital_signal_tr m_trans;

  	function new(string name, uvm_component parent);
  		super.new(name, parent);
  		analysis_port = new("analysis_port", this);
	endfunction
		
	// Methods run_phase, and do_mon generated by setting monitor_inc in file spi.tpl
	task run_phase(uvm_phase phase);
		`uvm_info(get_type_name(), "run_phase", UVM_HIGH)
		m_trans = digital_signal_tr::type_id::create("m_trans");
		do_mon();
	endtask
	
	`include "includes/digital_signal_monitor_inc.sv"
	
	// You can insert code here by setting monitor_inc_inside_class in file digital_signal.tpl
	
endclass

// You can insert code here by setting monitor_inc_after_class in file digital_signal.tpl

`endif

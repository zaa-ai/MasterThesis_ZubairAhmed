import buffer_if_pkg::*;
`include "DW_ecc_function.inc"

/**
 * Interface: clk_osc_if
 */
interface clk_osc_if;
	
	logic clk;
	
endinterface



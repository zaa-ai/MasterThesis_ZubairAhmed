/* ###   interface instances   ###################################################### */

TEST_OSC_TMR_ANA_TB_PLL_if TEST_OSC_TMR_ANA_TB_PLL (); 
TEST_OSC_TMR_ANA_TB_OSC_if TEST_OSC_TMR_ANA_TB_OSC (); 
TEST_OSC_TMR_DIG_TB_if TEST_OSC_TMR_DIG_TB (); 
TEST_OSC_TMR_VAL_TB_if TEST_OSC_TMR_VAL_TB (); 
TEST_OSC_TMR_SEL_TB_if TEST_OSC_TMR_SEL_TB (); 


typedef enum {L=0, H=1, X, Z} digital_signal_t ;


slave_timing[3][192+0].info_corner          = 3;
slave_timing[3][192+0].info_temp__j__       = -40;
slave_timing[3][192+0].info_i__quite_rec__  = 0.006000000;
slave_timing[3][192+0].info_dtr__ib__       = -1;
slave_timing[3][192+0].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+0].info_i__max_slave__  = 0.023000000;
slave_timing[3][192+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][192+0].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+0].t_rxd1[0][1] = 2728ns;
slave_timing[3][192+0].t_rxd1[1][0] = 2750ns;
slave_timing[3][192+0].t_rxd1[0][2] = 2044ns;
slave_timing[3][192+0].t_rxd1[2][0] = 3347ns;
slave_timing[3][192+0].t_rxd2[0][2] = 3296ns;
slave_timing[3][192+0].t_rxd2[2][0] = 2061ns;
slave_timing[3][192+0].t_rxd2[1][2] = 2686ns;
slave_timing[3][192+0].t_rxd2[2][1] = 2762ns;

slave_timing[3][192+1].info_corner          = 3;
slave_timing[3][192+1].info_temp__j__       = -40;
slave_timing[3][192+1].info_i__quite_rec__  = 0.006000000;
slave_timing[3][192+1].info_dtr__ib__       = -1;
slave_timing[3][192+1].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+1].info_i__max_slave__  = 0.025000000;
slave_timing[3][192+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][192+1].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+1].t_rxd1[0][1] = 2625ns;
slave_timing[3][192+1].t_rxd1[1][0] = 2837ns;
slave_timing[3][192+1].t_rxd1[0][2] = 1978ns;
slave_timing[3][192+1].t_rxd1[2][0] = 3408ns;
slave_timing[3][192+1].t_rxd2[0][2] = 3109ns;
slave_timing[3][192+1].t_rxd2[2][0] = 2210ns;
slave_timing[3][192+1].t_rxd2[1][2] = 2403ns;
slave_timing[3][192+1].t_rxd2[2][1] = 3004ns;

slave_timing[3][192+2].info_corner          = 3;
slave_timing[3][192+2].info_temp__j__       = -40;
slave_timing[3][192+2].info_i__quite_rec__  = 0.006000000;
slave_timing[3][192+2].info_dtr__ib__       = 1;
slave_timing[3][192+2].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+2].info_i__max_slave__  = 0.023000000;
slave_timing[3][192+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][192+2].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+2].t_rxd1[0][1] = 2812ns;
slave_timing[3][192+2].t_rxd1[1][0] = 2685ns;
slave_timing[3][192+2].t_rxd1[0][2] = 2088ns;
slave_timing[3][192+2].t_rxd1[2][0] = 3307ns;
slave_timing[3][192+2].t_rxd2[0][2] = 3467ns;
slave_timing[3][192+2].t_rxd2[2][0] = 1934ns;
slave_timing[3][192+2].t_rxd2[1][2] = 2933ns;
slave_timing[3][192+2].t_rxd2[2][1] = 2545ns;

slave_timing[3][192+3].info_corner          = 3;
slave_timing[3][192+3].info_temp__j__       = -40;
slave_timing[3][192+3].info_i__quite_rec__  = 0.006000000;
slave_timing[3][192+3].info_dtr__ib__       = 1;
slave_timing[3][192+3].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+3].info_i__max_slave__  = 0.025000000;
slave_timing[3][192+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][192+3].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+3].t_rxd1[0][1] = 2699ns;
slave_timing[3][192+3].t_rxd1[1][0] = 2773ns;
slave_timing[3][192+3].t_rxd1[0][2] = 2022ns;
slave_timing[3][192+3].t_rxd1[2][0] = 3363ns;
slave_timing[3][192+3].t_rxd2[0][2] = 3243ns;
slave_timing[3][192+3].t_rxd2[2][0] = 2103ns;
slave_timing[3][192+3].t_rxd2[1][2] = 2649ns;
slave_timing[3][192+3].t_rxd2[2][1] = 2792ns;

slave_timing[3][192+4].info_corner          = 3;
slave_timing[3][192+4].info_temp__j__       = -40;
slave_timing[3][192+4].info_i__quite_rec__  = 0.006000000;
slave_timing[3][192+4].info_dtr__ib__       = -1;
slave_timing[3][192+4].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+4].info_i__max_slave__  = 0.023000000;
slave_timing[3][192+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][192+4].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+4].t_rxd1[0][1] = 2808ns;
slave_timing[3][192+4].t_rxd1[1][0] = 2827ns;
slave_timing[3][192+4].t_rxd1[0][2] = 2115ns;
slave_timing[3][192+4].t_rxd1[2][0] = 3423ns;
slave_timing[3][192+4].t_rxd2[0][2] = 3311ns;
slave_timing[3][192+4].t_rxd2[2][0] = 2080ns;
slave_timing[3][192+4].t_rxd2[1][2] = 2703ns;
slave_timing[3][192+4].t_rxd2[2][1] = 2777ns;

slave_timing[3][192+5].info_corner          = 3;
slave_timing[3][192+5].info_temp__j__       = -40;
slave_timing[3][192+5].info_i__quite_rec__  = 0.006000000;
slave_timing[3][192+5].info_dtr__ib__       = -1;
slave_timing[3][192+5].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+5].info_i__max_slave__  = 0.025000000;
slave_timing[3][192+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][192+5].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+5].t_rxd1[0][1] = 2698ns;
slave_timing[3][192+5].t_rxd1[1][0] = 2909ns;
slave_timing[3][192+5].t_rxd1[0][2] = 2052ns;
slave_timing[3][192+5].t_rxd1[2][0] = 3480ns;
slave_timing[3][192+5].t_rxd2[0][2] = 3127ns;
slave_timing[3][192+5].t_rxd2[2][0] = 2224ns;
slave_timing[3][192+5].t_rxd2[1][2] = 2413ns;
slave_timing[3][192+5].t_rxd2[2][1] = 3063ns;

slave_timing[3][192+6].info_corner          = 3;
slave_timing[3][192+6].info_temp__j__       = -40;
slave_timing[3][192+6].info_i__quite_rec__  = 0.006000000;
slave_timing[3][192+6].info_dtr__ib__       = 1;
slave_timing[3][192+6].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+6].info_i__max_slave__  = 0.023000000;
slave_timing[3][192+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][192+6].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+6].t_rxd1[0][1] = 2880ns;
slave_timing[3][192+6].t_rxd1[1][0] = 2758ns;
slave_timing[3][192+6].t_rxd1[0][2] = 2152ns;
slave_timing[3][192+6].t_rxd1[2][0] = 3377ns;
slave_timing[3][192+6].t_rxd2[0][2] = 3479ns;
slave_timing[3][192+6].t_rxd2[2][0] = 1948ns;
slave_timing[3][192+6].t_rxd2[1][2] = 2984ns;
slave_timing[3][192+6].t_rxd2[2][1] = 2518ns;

slave_timing[3][192+7].info_corner          = 3;
slave_timing[3][192+7].info_temp__j__       = -40;
slave_timing[3][192+7].info_i__quite_rec__  = 0.006000000;
slave_timing[3][192+7].info_dtr__ib__       = 1;
slave_timing[3][192+7].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+7].info_i__max_slave__  = 0.025000000;
slave_timing[3][192+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][192+7].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+7].t_rxd1[0][1] = 2768ns;
slave_timing[3][192+7].t_rxd1[1][0] = 2844ns;
slave_timing[3][192+7].t_rxd1[0][2] = 2086ns;
slave_timing[3][192+7].t_rxd1[2][0] = 3431ns;
slave_timing[3][192+7].t_rxd2[0][2] = 3259ns;
slave_timing[3][192+7].t_rxd2[2][0] = 2113ns;
slave_timing[3][192+7].t_rxd2[1][2] = 2619ns;
slave_timing[3][192+7].t_rxd2[2][1] = 2846ns;

slave_timing[3][192+8].info_corner          = 3;
slave_timing[3][192+8].info_temp__j__       = -40;
slave_timing[3][192+8].info_i__quite_rec__  = 0.003000000;
slave_timing[3][192+8].info_dtr__ib__       = -1;
slave_timing[3][192+8].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+8].info_i__max_slave__  = 0.023000000;
slave_timing[3][192+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][192+8].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+8].t_rxd1[0][1] = 2755ns;
slave_timing[3][192+8].t_rxd1[1][0] = 2727ns;
slave_timing[3][192+8].t_rxd1[0][2] = 2039ns;
slave_timing[3][192+8].t_rxd1[2][0] = 3359ns;
slave_timing[3][192+8].t_rxd2[0][2] = 3292ns;
slave_timing[3][192+8].t_rxd2[2][0] = 2071ns;
slave_timing[3][192+8].t_rxd2[1][2] = 2719ns;
slave_timing[3][192+8].t_rxd2[2][1] = 2732ns;

slave_timing[3][192+9].info_corner          = 3;
slave_timing[3][192+9].info_temp__j__       = -40;
slave_timing[3][192+9].info_i__quite_rec__  = 0.003000000;
slave_timing[3][192+9].info_dtr__ib__       = -1;
slave_timing[3][192+9].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+9].info_i__max_slave__  = 0.025000000;
slave_timing[3][192+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][192+9].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+9].t_rxd1[0][1] = 2617ns;
slave_timing[3][192+9].t_rxd1[1][0] = 2848ns;
slave_timing[3][192+9].t_rxd1[0][2] = 1975ns;
slave_timing[3][192+9].t_rxd1[2][0] = 3413ns;
slave_timing[3][192+9].t_rxd2[0][2] = 3104ns;
slave_timing[3][192+9].t_rxd2[2][0] = 2210ns;
slave_timing[3][192+9].t_rxd2[1][2] = 2391ns;
slave_timing[3][192+9].t_rxd2[2][1] = 3055ns;

slave_timing[3][192+10].info_corner          = 3;
slave_timing[3][192+10].info_temp__j__       = -40;
slave_timing[3][192+10].info_i__quite_rec__  = 0.003000000;
slave_timing[3][192+10].info_dtr__ib__       = 1;
slave_timing[3][192+10].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+10].info_i__max_slave__  = 0.023000000;
slave_timing[3][192+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][192+10].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+10].t_rxd1[0][1] = 2795ns;
slave_timing[3][192+10].t_rxd1[1][0] = 2692ns;
slave_timing[3][192+10].t_rxd1[0][2] = 2082ns;
slave_timing[3][192+10].t_rxd1[2][0] = 3319ns;
slave_timing[3][192+10].t_rxd2[0][2] = 3453ns;
slave_timing[3][192+10].t_rxd2[2][0] = 1941ns;
slave_timing[3][192+10].t_rxd2[1][2] = 2924ns;
slave_timing[3][192+10].t_rxd2[2][1] = 2552ns;

slave_timing[3][192+11].info_corner          = 3;
slave_timing[3][192+11].info_temp__j__       = -40;
slave_timing[3][192+11].info_i__quite_rec__  = 0.003000000;
slave_timing[3][192+11].info_dtr__ib__       = 1;
slave_timing[3][192+11].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+11].info_i__max_slave__  = 0.025000000;
slave_timing[3][192+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][192+11].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+11].t_rxd1[0][1] = 2689ns;
slave_timing[3][192+11].t_rxd1[1][0] = 2780ns;
slave_timing[3][192+11].t_rxd1[0][2] = 2014ns;
slave_timing[3][192+11].t_rxd1[2][0] = 3368ns;
slave_timing[3][192+11].t_rxd2[0][2] = 3234ns;
slave_timing[3][192+11].t_rxd2[2][0] = 2107ns;
slave_timing[3][192+11].t_rxd2[1][2] = 2601ns;
slave_timing[3][192+11].t_rxd2[2][1] = 2839ns;

slave_timing[3][192+12].info_corner          = 3;
slave_timing[3][192+12].info_temp__j__       = -40;
slave_timing[3][192+12].info_i__quite_rec__  = 0.003000000;
slave_timing[3][192+12].info_dtr__ib__       = -1;
slave_timing[3][192+12].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+12].info_i__max_slave__  = 0.023000000;
slave_timing[3][192+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][192+12].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+12].t_rxd1[0][1] = 2799ns;
slave_timing[3][192+12].t_rxd1[1][0] = 2844ns;
slave_timing[3][192+12].t_rxd1[0][2] = 2116ns;
slave_timing[3][192+12].t_rxd1[2][0] = 3437ns;
slave_timing[3][192+12].t_rxd2[0][2] = 3304ns;
slave_timing[3][192+12].t_rxd2[2][0] = 2083ns;
slave_timing[3][192+12].t_rxd2[1][2] = 2730ns;
slave_timing[3][192+12].t_rxd2[2][1] = 2739ns;

slave_timing[3][192+13].info_corner          = 3;
slave_timing[3][192+13].info_temp__j__       = -40;
slave_timing[3][192+13].info_i__quite_rec__  = 0.003000000;
slave_timing[3][192+13].info_dtr__ib__       = -1;
slave_timing[3][192+13].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+13].info_i__max_slave__  = 0.025000000;
slave_timing[3][192+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][192+13].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+13].t_rxd1[0][1] = 2693ns;
slave_timing[3][192+13].t_rxd1[1][0] = 2924ns;
slave_timing[3][192+13].t_rxd1[0][2] = 2049ns;
slave_timing[3][192+13].t_rxd1[2][0] = 3492ns;
slave_timing[3][192+13].t_rxd2[0][2] = 3117ns;
slave_timing[3][192+13].t_rxd2[2][0] = 2229ns;
slave_timing[3][192+13].t_rxd2[1][2] = 2408ns;
slave_timing[3][192+13].t_rxd2[2][1] = 3070ns;

slave_timing[3][192+14].info_corner          = 3;
slave_timing[3][192+14].info_temp__j__       = -40;
slave_timing[3][192+14].info_i__quite_rec__  = 0.003000000;
slave_timing[3][192+14].info_dtr__ib__       = 1;
slave_timing[3][192+14].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+14].info_i__max_slave__  = 0.023000000;
slave_timing[3][192+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][192+14].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+14].t_rxd1[0][1] = 2871ns;
slave_timing[3][192+14].t_rxd1[1][0] = 2757ns;
slave_timing[3][192+14].t_rxd1[0][2] = 2154ns;
slave_timing[3][192+14].t_rxd1[2][0] = 3380ns;
slave_timing[3][192+14].t_rxd2[0][2] = 3467ns;
slave_timing[3][192+14].t_rxd2[2][0] = 1954ns;
slave_timing[3][192+14].t_rxd2[1][2] = 2975ns;
slave_timing[3][192+14].t_rxd2[2][1] = 2526ns;

slave_timing[3][192+15].info_corner          = 3;
slave_timing[3][192+15].info_temp__j__       = -40;
slave_timing[3][192+15].info_i__quite_rec__  = 0.003000000;
slave_timing[3][192+15].info_dtr__ib__       = 1;
slave_timing[3][192+15].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+15].info_i__max_slave__  = 0.025000000;
slave_timing[3][192+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][192+15].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+15].t_rxd1[0][1] = 2799ns;
slave_timing[3][192+15].t_rxd1[1][0] = 2811ns;
slave_timing[3][192+15].t_rxd1[0][2] = 2085ns;
slave_timing[3][192+15].t_rxd1[2][0] = 3438ns;
slave_timing[3][192+15].t_rxd2[0][2] = 3251ns;
slave_timing[3][192+15].t_rxd2[2][0] = 2121ns;
slave_timing[3][192+15].t_rxd2[1][2] = 2652ns;
slave_timing[3][192+15].t_rxd2[2][1] = 2812ns;

slave_timing[3][192+16].info_corner          = 3;
slave_timing[3][192+16].info_temp__j__       = -40;
slave_timing[3][192+16].info_i__quite_rec__  = 0.000000000;
slave_timing[3][192+16].info_dtr__ib__       = -1;
slave_timing[3][192+16].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+16].info_i__max_slave__  = 0.023000000;
slave_timing[3][192+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][192+16].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+16].t_rxd1[0][1] = 2743ns;
slave_timing[3][192+16].t_rxd1[1][0] = 2737ns;
slave_timing[3][192+16].t_rxd1[0][2] = 2051ns;
slave_timing[3][192+16].t_rxd1[2][0] = 3339ns;
slave_timing[3][192+16].t_rxd2[0][2] = 3306ns;
slave_timing[3][192+16].t_rxd2[2][0] = 2056ns;
slave_timing[3][192+16].t_rxd2[1][2] = 2707ns;
slave_timing[3][192+16].t_rxd2[2][1] = 2742ns;

slave_timing[3][192+17].info_corner          = 3;
slave_timing[3][192+17].info_temp__j__       = -40;
slave_timing[3][192+17].info_i__quite_rec__  = 0.000000000;
slave_timing[3][192+17].info_dtr__ib__       = -1;
slave_timing[3][192+17].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+17].info_i__max_slave__  = 0.025000000;
slave_timing[3][192+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][192+17].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+17].t_rxd1[0][1] = 2636ns;
slave_timing[3][192+17].t_rxd1[1][0] = 2815ns;
slave_timing[3][192+17].t_rxd1[0][2] = 1989ns;
slave_timing[3][192+17].t_rxd1[2][0] = 3396ns;
slave_timing[3][192+17].t_rxd2[0][2] = 3119ns;
slave_timing[3][192+17].t_rxd2[2][0] = 2201ns;
slave_timing[3][192+17].t_rxd2[1][2] = 2415ns;
slave_timing[3][192+17].t_rxd2[2][1] = 3032ns;

slave_timing[3][192+18].info_corner          = 3;
slave_timing[3][192+18].info_temp__j__       = -40;
slave_timing[3][192+18].info_i__quite_rec__  = 0.000000000;
slave_timing[3][192+18].info_dtr__ib__       = 1;
slave_timing[3][192+18].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+18].info_i__max_slave__  = 0.023000000;
slave_timing[3][192+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][192+18].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+18].t_rxd1[0][1] = 2831ns;
slave_timing[3][192+18].t_rxd1[1][0] = 2664ns;
slave_timing[3][192+18].t_rxd1[0][2] = 2099ns;
slave_timing[3][192+18].t_rxd1[2][0] = 3295ns;
slave_timing[3][192+18].t_rxd2[0][2] = 3477ns;
slave_timing[3][192+18].t_rxd2[2][0] = 1920ns;
slave_timing[3][192+18].t_rxd2[1][2] = 2957ns;
slave_timing[3][192+18].t_rxd2[2][1] = 2477ns;

slave_timing[3][192+19].info_corner          = 3;
slave_timing[3][192+19].info_temp__j__       = -40;
slave_timing[3][192+19].info_i__quite_rec__  = 0.000000000;
slave_timing[3][192+19].info_dtr__ib__       = 1;
slave_timing[3][192+19].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+19].info_i__max_slave__  = 0.025000000;
slave_timing[3][192+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][192+19].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+19].t_rxd1[0][1] = 2716ns;
slave_timing[3][192+19].t_rxd1[1][0] = 2752ns;
slave_timing[3][192+19].t_rxd1[0][2] = 2035ns;
slave_timing[3][192+19].t_rxd1[2][0] = 3350ns;
slave_timing[3][192+19].t_rxd2[0][2] = 3253ns;
slave_timing[3][192+19].t_rxd2[2][0] = 2088ns;
slave_timing[3][192+19].t_rxd2[1][2] = 2626ns;
slave_timing[3][192+19].t_rxd2[2][1] = 2807ns;

slave_timing[3][192+20].info_corner          = 3;
slave_timing[3][192+20].info_temp__j__       = -40;
slave_timing[3][192+20].info_i__quite_rec__  = 0.000000000;
slave_timing[3][192+20].info_dtr__ib__       = -1;
slave_timing[3][192+20].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+20].info_i__max_slave__  = 0.023000000;
slave_timing[3][192+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][192+20].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+20].t_rxd1[0][1] = 2827ns;
slave_timing[3][192+20].t_rxd1[1][0] = 2810ns;
slave_timing[3][192+20].t_rxd1[0][2] = 2126ns;
slave_timing[3][192+20].t_rxd1[2][0] = 3410ns;
slave_timing[3][192+20].t_rxd2[0][2] = 3317ns;
slave_timing[3][192+20].t_rxd2[2][0] = 2071ns;
slave_timing[3][192+20].t_rxd2[1][2] = 2717ns;
slave_timing[3][192+20].t_rxd2[2][1] = 2749ns;

slave_timing[3][192+21].info_corner          = 3;
slave_timing[3][192+21].info_temp__j__       = -40;
slave_timing[3][192+21].info_i__quite_rec__  = 0.000000000;
slave_timing[3][192+21].info_dtr__ib__       = -1;
slave_timing[3][192+21].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+21].info_i__max_slave__  = 0.025000000;
slave_timing[3][192+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][192+21].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+21].t_rxd1[0][1] = 2719ns;
slave_timing[3][192+21].t_rxd1[1][0] = 2892ns;
slave_timing[3][192+21].t_rxd1[0][2] = 2065ns;
slave_timing[3][192+21].t_rxd1[2][0] = 3471ns;
slave_timing[3][192+21].t_rxd2[0][2] = 3131ns;
slave_timing[3][192+21].t_rxd2[2][0] = 2211ns;
slave_timing[3][192+21].t_rxd2[1][2] = 2430ns;
slave_timing[3][192+21].t_rxd2[2][1] = 3000ns;

slave_timing[3][192+22].info_corner          = 3;
slave_timing[3][192+22].info_temp__j__       = -40;
slave_timing[3][192+22].info_i__quite_rec__  = 0.000000000;
slave_timing[3][192+22].info_dtr__ib__       = 1;
slave_timing[3][192+22].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+22].info_i__max_slave__  = 0.023000000;
slave_timing[3][192+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][192+22].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+22].t_rxd1[0][1] = 2901ns;
slave_timing[3][192+22].t_rxd1[1][0] = 2736ns;
slave_timing[3][192+22].t_rxd1[0][2] = 2166ns;
slave_timing[3][192+22].t_rxd1[2][0] = 3361ns;
slave_timing[3][192+22].t_rxd2[0][2] = 3487ns;
slave_timing[3][192+22].t_rxd2[2][0] = 1932ns;
slave_timing[3][192+22].t_rxd2[1][2] = 3014ns;
slave_timing[3][192+22].t_rxd2[2][1] = 2496ns;

slave_timing[3][192+23].info_corner          = 3;
slave_timing[3][192+23].info_temp__j__       = -40;
slave_timing[3][192+23].info_i__quite_rec__  = 0.000000000;
slave_timing[3][192+23].info_dtr__ib__       = 1;
slave_timing[3][192+23].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+23].info_i__max_slave__  = 0.025000000;
slave_timing[3][192+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][192+23].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+23].t_rxd1[0][1] = 2788ns;
slave_timing[3][192+23].t_rxd1[1][0] = 2821ns;
slave_timing[3][192+23].t_rxd1[0][2] = 2102ns;
slave_timing[3][192+23].t_rxd1[2][0] = 3419ns;
slave_timing[3][192+23].t_rxd2[0][2] = 3267ns;
slave_timing[3][192+23].t_rxd2[2][0] = 2098ns;
slave_timing[3][192+23].t_rxd2[1][2] = 2640ns;
slave_timing[3][192+23].t_rxd2[2][1] = 2821ns;

slave_timing[3][192+24].info_corner          = 3;
slave_timing[3][192+24].info_temp__j__       = -40;
slave_timing[3][192+24].info_i__quite_rec__  = 0.040000000;
slave_timing[3][192+24].info_dtr__ib__       = -1;
slave_timing[3][192+24].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+24].info_i__max_slave__  = 0.023000000;
slave_timing[3][192+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][192+24].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+24].t_rxd1[0][1] = 2740ns;
slave_timing[3][192+24].t_rxd1[1][0] = 2717ns;
slave_timing[3][192+24].t_rxd1[0][2] = 2048ns;
slave_timing[3][192+24].t_rxd1[2][0] = 3322ns;
slave_timing[3][192+24].t_rxd2[0][2] = 3310ns;
slave_timing[3][192+24].t_rxd2[2][0] = 2050ns;
slave_timing[3][192+24].t_rxd2[1][2] = 2713ns;
slave_timing[3][192+24].t_rxd2[2][1] = 2730ns;

slave_timing[3][192+25].info_corner          = 3;
slave_timing[3][192+25].info_temp__j__       = -40;
slave_timing[3][192+25].info_i__quite_rec__  = 0.040000000;
slave_timing[3][192+25].info_dtr__ib__       = -1;
slave_timing[3][192+25].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+25].info_i__max_slave__  = 0.025000000;
slave_timing[3][192+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][192+25].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+25].t_rxd1[0][1] = 2637ns;
slave_timing[3][192+25].t_rxd1[1][0] = 2800ns;
slave_timing[3][192+25].t_rxd1[0][2] = 1983ns;
slave_timing[3][192+25].t_rxd1[2][0] = 3376ns;
slave_timing[3][192+25].t_rxd2[0][2] = 3124ns;
slave_timing[3][192+25].t_rxd2[2][0] = 2196ns;
slave_timing[3][192+25].t_rxd2[1][2] = 2428ns;
slave_timing[3][192+25].t_rxd2[2][1] = 2981ns;

slave_timing[3][192+26].info_corner          = 3;
slave_timing[3][192+26].info_temp__j__       = -40;
slave_timing[3][192+26].info_i__quite_rec__  = 0.040000000;
slave_timing[3][192+26].info_dtr__ib__       = 1;
slave_timing[3][192+26].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+26].info_i__max_slave__  = 0.023000000;
slave_timing[3][192+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][192+26].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+26].t_rxd1[0][1] = 2817ns;
slave_timing[3][192+26].t_rxd1[1][0] = 2659ns;
slave_timing[3][192+26].t_rxd1[0][2] = 2089ns;
slave_timing[3][192+26].t_rxd1[2][0] = 3286ns;
slave_timing[3][192+26].t_rxd2[0][2] = 3477ns;
slave_timing[3][192+26].t_rxd2[2][0] = 1923ns;
slave_timing[3][192+26].t_rxd2[1][2] = 2955ns;
slave_timing[3][192+26].t_rxd2[2][1] = 2520ns;

slave_timing[3][192+27].info_corner          = 3;
slave_timing[3][192+27].info_temp__j__       = -40;
slave_timing[3][192+27].info_i__quite_rec__  = 0.040000000;
slave_timing[3][192+27].info_dtr__ib__       = 1;
slave_timing[3][192+27].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+27].info_i__max_slave__  = 0.025000000;
slave_timing[3][192+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[3][192+27].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+27].t_rxd1[0][1] = 2705ns;
slave_timing[3][192+27].t_rxd1[1][0] = 2748ns;
slave_timing[3][192+27].t_rxd1[0][2] = 2025ns;
slave_timing[3][192+27].t_rxd1[2][0] = 3344ns;
slave_timing[3][192+27].t_rxd2[0][2] = 3253ns;
slave_timing[3][192+27].t_rxd2[2][0] = 2092ns;
slave_timing[3][192+27].t_rxd2[1][2] = 2629ns;
slave_timing[3][192+27].t_rxd2[2][1] = 2815ns;

slave_timing[3][192+28].info_corner          = 3;
slave_timing[3][192+28].info_temp__j__       = -40;
slave_timing[3][192+28].info_i__quite_rec__  = 0.040000000;
slave_timing[3][192+28].info_dtr__ib__       = -1;
slave_timing[3][192+28].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+28].info_i__max_slave__  = 0.023000000;
slave_timing[3][192+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][192+28].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+28].t_rxd1[0][1] = 2790ns;
slave_timing[3][192+28].t_rxd1[1][0] = 2763ns;
slave_timing[3][192+28].t_rxd1[0][2] = 2088ns;
slave_timing[3][192+28].t_rxd1[2][0] = 3366ns;
slave_timing[3][192+28].t_rxd2[0][2] = 3324ns;
slave_timing[3][192+28].t_rxd2[2][0] = 2063ns;
slave_timing[3][192+28].t_rxd2[1][2] = 2731ns;
slave_timing[3][192+28].t_rxd2[2][1] = 2744ns;

slave_timing[3][192+29].info_corner          = 3;
slave_timing[3][192+29].info_temp__j__       = -40;
slave_timing[3][192+29].info_i__quite_rec__  = 0.040000000;
slave_timing[3][192+29].info_dtr__ib__       = -1;
slave_timing[3][192+29].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+29].info_i__max_slave__  = 0.025000000;
slave_timing[3][192+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][192+29].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+29].t_rxd1[0][1] = 2684ns;
slave_timing[3][192+29].t_rxd1[1][0] = 2843ns;
slave_timing[3][192+29].t_rxd1[0][2] = 2022ns;
slave_timing[3][192+29].t_rxd1[2][0] = 3423ns;
slave_timing[3][192+29].t_rxd2[0][2] = 3139ns;
slave_timing[3][192+29].t_rxd2[2][0] = 2210ns;
slave_timing[3][192+29].t_rxd2[1][2] = 2439ns;
slave_timing[3][192+29].t_rxd2[2][1] = 3034ns;

slave_timing[3][192+30].info_corner          = 3;
slave_timing[3][192+30].info_temp__j__       = -40;
slave_timing[3][192+30].info_i__quite_rec__  = 0.040000000;
slave_timing[3][192+30].info_dtr__ib__       = 1;
slave_timing[3][192+30].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+30].info_i__max_slave__  = 0.023000000;
slave_timing[3][192+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][192+30].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+30].t_rxd1[0][1] = 2860ns;
slave_timing[3][192+30].t_rxd1[1][0] = 2701ns;
slave_timing[3][192+30].t_rxd1[0][2] = 2126ns;
slave_timing[3][192+30].t_rxd1[2][0] = 3328ns;
slave_timing[3][192+30].t_rxd2[0][2] = 3490ns;
slave_timing[3][192+30].t_rxd2[2][0] = 1932ns;
slave_timing[3][192+30].t_rxd2[1][2] = 2966ns;
slave_timing[3][192+30].t_rxd2[2][1] = 2540ns;

slave_timing[3][192+31].info_corner          = 3;
slave_timing[3][192+31].info_temp__j__       = -40;
slave_timing[3][192+31].info_i__quite_rec__  = 0.040000000;
slave_timing[3][192+31].info_dtr__ib__       = 1;
slave_timing[3][192+31].info_i__offset_rec__ = 0.000000000;
slave_timing[3][192+31].info_i__max_slave__  = 0.025000000;
slave_timing[3][192+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[3][192+31].info_r__dsi_bus__    = 5.000;

slave_timing[3][192+31].t_rxd1[0][1] = 2746ns;
slave_timing[3][192+31].t_rxd1[1][0] = 2787ns;
slave_timing[3][192+31].t_rxd1[0][2] = 2062ns;
slave_timing[3][192+31].t_rxd1[2][0] = 3382ns;
slave_timing[3][192+31].t_rxd2[0][2] = 3267ns;
slave_timing[3][192+31].t_rxd2[2][0] = 2103ns;
slave_timing[3][192+31].t_rxd2[1][2] = 2640ns;
slave_timing[3][192+31].t_rxd2[2][1] = 2825ns;

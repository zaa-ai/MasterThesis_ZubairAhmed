/* ###   interface instances   ###################################################### */

DSI3_channel_trimming_registers_TRIM_DSI_REC_FALL_if DSI3_channel_trimming_registers_TRIM_DSI_REC_FALL (); 
DSI3_channel_trimming_registers_TRIM_DSI_REC_RISE_if DSI3_channel_trimming_registers_TRIM_DSI_REC_RISE (); 


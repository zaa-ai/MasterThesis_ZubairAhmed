/* ###   interface instances   ###################################################### */

IC_revision_and_ID_registers_CHIP_ID_LOW_if IC_revision_and_ID_registers_CHIP_ID_LOW (); 
IC_revision_and_ID_registers_CHIP_ID_HIGH_if IC_revision_and_ID_registers_CHIP_ID_HIGH (); 
IC_revision_and_ID_registers_IC_REVISION_if IC_revision_and_ID_registers_IC_REVISION (); 


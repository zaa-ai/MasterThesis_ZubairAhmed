/* ###   interface instances   ###################################################### */

DSI3_channel_registers_DSI_STAT_if DSI3_channel_registers_DSI_STAT (); 
DSI3_channel_registers_PDCM_PERIOD_if DSI3_channel_registers_PDCM_PERIOD (); 
DSI3_channel_registers_DSI_LOAD_if DSI3_channel_registers_DSI_LOAD (); 
DSI3_channel_registers_DSI_IRQ_STAT_if DSI3_channel_registers_DSI_IRQ_STAT (); 
DSI3_channel_registers_DSI_IRQ_MASK_if DSI3_channel_registers_DSI_IRQ_MASK (); 
DSI3_channel_registers_DSI_CMD_if DSI3_channel_registers_DSI_CMD (); 
DSI3_channel_registers_CRM_WORD2_if DSI3_channel_registers_CRM_WORD2 (); 
DSI3_channel_registers_CRM_WORD1_if DSI3_channel_registers_CRM_WORD1 (); 
DSI3_channel_registers_PACKET_STAT_if DSI3_channel_registers_PACKET_STAT (); 
DSI3_channel_registers_WAIT_TIME_if DSI3_channel_registers_WAIT_TIME (); 
DSI3_channel_registers_SYNC_if DSI3_channel_registers_SYNC (); 
DSI3_channel_registers_FRAME_STAT_if DSI3_channel_registers_FRAME_STAT (); 


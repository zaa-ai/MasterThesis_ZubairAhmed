/* ###   interface instances   ###################################################### */

SPI_registers_SPI_IRQ_STAT_if SPI_registers_SPI_IRQ_STAT (); 
SPI_registers_SPI_IRQ_MASK_if SPI_registers_SPI_IRQ_MASK (); 
SPI_registers_STATUS_WORD_if SPI_registers_STATUS_WORD (); 


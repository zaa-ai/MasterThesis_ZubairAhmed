/**
 * Interface: OTP_model_if
 * 
 * TODO: Add interface documentation
 */
interface OTP_model_if;

	string dat_file;
	
endinterface



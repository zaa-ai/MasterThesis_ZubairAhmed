
slave_timing[0][160+0].info_corner          = 2;
slave_timing[0][160+0].info_temp__j__       = -40;
slave_timing[0][160+0].info_i__quite_rec__  = 0.006000000;
slave_timing[0][160+0].info_dtr__ib__       = -1;
slave_timing[0][160+0].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+0].info_i__max_slave__  = 0.023000000;
slave_timing[0][160+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][160+0].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+0].t_rxd1[0][1] = 1097ns;
slave_timing[0][160+0].t_rxd1[1][0] = 1111ns;
slave_timing[0][160+0].t_rxd1[0][2] = 807ns;
slave_timing[0][160+0].t_rxd1[2][0] = 1401ns;
slave_timing[0][160+0].t_rxd2[0][2] = 1363ns;
slave_timing[0][160+0].t_rxd2[2][0] = 815ns;
slave_timing[0][160+0].t_rxd2[1][2] = 1077ns;
slave_timing[0][160+0].t_rxd2[2][1] = 1100ns;

slave_timing[0][160+1].info_corner          = 2;
slave_timing[0][160+1].info_temp__j__       = -40;
slave_timing[0][160+1].info_i__quite_rec__  = 0.006000000;
slave_timing[0][160+1].info_dtr__ib__       = -1;
slave_timing[0][160+1].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+1].info_i__max_slave__  = 0.025000000;
slave_timing[0][160+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][160+1].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+1].t_rxd1[0][1] = 1050ns;
slave_timing[0][160+1].t_rxd1[1][0] = 1150ns;
slave_timing[0][160+1].t_rxd1[0][2] = 785ns;
slave_timing[0][160+1].t_rxd1[2][0] = 1432ns;
slave_timing[0][160+1].t_rxd2[0][2] = 1263ns;
slave_timing[0][160+1].t_rxd2[2][0] = 870ns;
slave_timing[0][160+1].t_rxd2[1][2] = 950ns;
slave_timing[0][160+1].t_rxd2[2][1] = 1233ns;

slave_timing[0][160+2].info_corner          = 2;
slave_timing[0][160+2].info_temp__j__       = -40;
slave_timing[0][160+2].info_i__quite_rec__  = 0.006000000;
slave_timing[0][160+2].info_dtr__ib__       = 1;
slave_timing[0][160+2].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+2].info_i__max_slave__  = 0.023000000;
slave_timing[0][160+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][160+2].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+2].t_rxd1[0][1] = 1133ns;
slave_timing[0][160+2].t_rxd1[1][0] = 1083ns;
slave_timing[0][160+2].t_rxd1[0][2] = 824ns;
slave_timing[0][160+2].t_rxd1[2][0] = 1377ns;
slave_timing[0][160+2].t_rxd2[0][2] = 1459ns;
slave_timing[0][160+2].t_rxd2[2][0] = 770ns;
slave_timing[0][160+2].t_rxd2[1][2] = 1190ns;
slave_timing[0][160+2].t_rxd2[2][1] = 1006ns;

slave_timing[0][160+3].info_corner          = 2;
slave_timing[0][160+3].info_temp__j__       = -40;
slave_timing[0][160+3].info_i__quite_rec__  = 0.006000000;
slave_timing[0][160+3].info_dtr__ib__       = 1;
slave_timing[0][160+3].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+3].info_i__max_slave__  = 0.025000000;
slave_timing[0][160+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][160+3].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+3].t_rxd1[0][1] = 1081ns;
slave_timing[0][160+3].t_rxd1[1][0] = 1121ns;
slave_timing[0][160+3].t_rxd1[0][2] = 798ns;
slave_timing[0][160+3].t_rxd1[2][0] = 1407ns;
slave_timing[0][160+3].t_rxd2[0][2] = 1332ns;
slave_timing[0][160+3].t_rxd2[2][0] = 830ns;
slave_timing[0][160+3].t_rxd2[1][2] = 1043ns;
slave_timing[0][160+3].t_rxd2[2][1] = 1132ns;

slave_timing[0][160+4].info_corner          = 2;
slave_timing[0][160+4].info_temp__j__       = -40;
slave_timing[0][160+4].info_i__quite_rec__  = 0.006000000;
slave_timing[0][160+4].info_dtr__ib__       = -1;
slave_timing[0][160+4].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+4].info_i__max_slave__  = 0.023000000;
slave_timing[0][160+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][160+4].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+4].t_rxd1[0][1] = 1169ns;
slave_timing[0][160+4].t_rxd1[1][0] = 1183ns;
slave_timing[0][160+4].t_rxd1[0][2] = 863ns;
slave_timing[0][160+4].t_rxd1[2][0] = 1462ns;
slave_timing[0][160+4].t_rxd2[0][2] = 1385ns;
slave_timing[0][160+4].t_rxd2[2][0] = 834ns;
slave_timing[0][160+4].t_rxd2[1][2] = 1089ns;
slave_timing[0][160+4].t_rxd2[2][1] = 1108ns;

slave_timing[0][160+5].info_corner          = 2;
slave_timing[0][160+5].info_temp__j__       = -40;
slave_timing[0][160+5].info_i__quite_rec__  = 0.006000000;
slave_timing[0][160+5].info_dtr__ib__       = -1;
slave_timing[0][160+5].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+5].info_i__max_slave__  = 0.025000000;
slave_timing[0][160+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][160+5].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+5].t_rxd1[0][1] = 1119ns;
slave_timing[0][160+5].t_rxd1[1][0] = 1220ns;
slave_timing[0][160+5].t_rxd1[0][2] = 838ns;
slave_timing[0][160+5].t_rxd1[2][0] = 1492ns;
slave_timing[0][160+5].t_rxd2[0][2] = 1286ns;
slave_timing[0][160+5].t_rxd2[2][0] = 887ns;
slave_timing[0][160+5].t_rxd2[1][2] = 966ns;
slave_timing[0][160+5].t_rxd2[2][1] = 1240ns;

slave_timing[0][160+6].info_corner          = 2;
slave_timing[0][160+6].info_temp__j__       = -40;
slave_timing[0][160+6].info_i__quite_rec__  = 0.006000000;
slave_timing[0][160+6].info_dtr__ib__       = 1;
slave_timing[0][160+6].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+6].info_i__max_slave__  = 0.023000000;
slave_timing[0][160+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][160+6].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+6].t_rxd1[0][1] = 1200ns;
slave_timing[0][160+6].t_rxd1[1][0] = 1148ns;
slave_timing[0][160+6].t_rxd1[0][2] = 874ns;
slave_timing[0][160+6].t_rxd1[2][0] = 1434ns;
slave_timing[0][160+6].t_rxd2[0][2] = 1477ns;
slave_timing[0][160+6].t_rxd2[2][0] = 785ns;
slave_timing[0][160+6].t_rxd2[1][2] = 1196ns;
slave_timing[0][160+6].t_rxd2[2][1] = 1019ns;

slave_timing[0][160+7].info_corner          = 2;
slave_timing[0][160+7].info_temp__j__       = -40;
slave_timing[0][160+7].info_i__quite_rec__  = 0.006000000;
slave_timing[0][160+7].info_dtr__ib__       = 1;
slave_timing[0][160+7].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+7].info_i__max_slave__  = 0.025000000;
slave_timing[0][160+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][160+7].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+7].t_rxd1[0][1] = 1145ns;
slave_timing[0][160+7].t_rxd1[1][0] = 1187ns;
slave_timing[0][160+7].t_rxd1[0][2] = 849ns;
slave_timing[0][160+7].t_rxd1[2][0] = 1464ns;
slave_timing[0][160+7].t_rxd2[0][2] = 1352ns;
slave_timing[0][160+7].t_rxd2[2][0] = 846ns;
slave_timing[0][160+7].t_rxd2[1][2] = 1052ns;
slave_timing[0][160+7].t_rxd2[2][1] = 1141ns;

slave_timing[0][160+8].info_corner          = 2;
slave_timing[0][160+8].info_temp__j__       = -40;
slave_timing[0][160+8].info_i__quite_rec__  = 0.003000000;
slave_timing[0][160+8].info_dtr__ib__       = -1;
slave_timing[0][160+8].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+8].info_i__max_slave__  = 0.023000000;
slave_timing[0][160+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][160+8].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+8].t_rxd1[0][1] = 1090ns;
slave_timing[0][160+8].t_rxd1[1][0] = 1119ns;
slave_timing[0][160+8].t_rxd1[0][2] = 804ns;
slave_timing[0][160+8].t_rxd1[2][0] = 1406ns;
slave_timing[0][160+8].t_rxd2[0][2] = 1358ns;
slave_timing[0][160+8].t_rxd2[2][0] = 821ns;
slave_timing[0][160+8].t_rxd2[1][2] = 1071ns;
slave_timing[0][160+8].t_rxd2[2][1] = 1109ns;

slave_timing[0][160+9].info_corner          = 2;
slave_timing[0][160+9].info_temp__j__       = -40;
slave_timing[0][160+9].info_i__quite_rec__  = 0.003000000;
slave_timing[0][160+9].info_dtr__ib__       = -1;
slave_timing[0][160+9].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+9].info_i__max_slave__  = 0.025000000;
slave_timing[0][160+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][160+9].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+9].t_rxd1[0][1] = 1041ns;
slave_timing[0][160+9].t_rxd1[1][0] = 1154ns;
slave_timing[0][160+9].t_rxd1[0][2] = 780ns;
slave_timing[0][160+9].t_rxd1[2][0] = 1436ns;
slave_timing[0][160+9].t_rxd2[0][2] = 1259ns;
slave_timing[0][160+9].t_rxd2[2][0] = 873ns;
slave_timing[0][160+9].t_rxd2[1][2] = 947ns;
slave_timing[0][160+9].t_rxd2[2][1] = 1247ns;

slave_timing[0][160+10].info_corner          = 2;
slave_timing[0][160+10].info_temp__j__       = -40;
slave_timing[0][160+10].info_i__quite_rec__  = 0.003000000;
slave_timing[0][160+10].info_dtr__ib__       = 1;
slave_timing[0][160+10].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+10].info_i__max_slave__  = 0.023000000;
slave_timing[0][160+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][160+10].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+10].t_rxd1[0][1] = 1124ns;
slave_timing[0][160+10].t_rxd1[1][0] = 1090ns;
slave_timing[0][160+10].t_rxd1[0][2] = 816ns;
slave_timing[0][160+10].t_rxd1[2][0] = 1381ns;
slave_timing[0][160+10].t_rxd2[0][2] = 1452ns;
slave_timing[0][160+10].t_rxd2[2][0] = 774ns;
slave_timing[0][160+10].t_rxd2[1][2] = 1181ns;
slave_timing[0][160+10].t_rxd2[2][1] = 1016ns;

slave_timing[0][160+11].info_corner          = 2;
slave_timing[0][160+11].info_temp__j__       = -40;
slave_timing[0][160+11].info_i__quite_rec__  = 0.003000000;
slave_timing[0][160+11].info_dtr__ib__       = 1;
slave_timing[0][160+11].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+11].info_i__max_slave__  = 0.025000000;
slave_timing[0][160+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][160+11].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+11].t_rxd1[0][1] = 1075ns;
slave_timing[0][160+11].t_rxd1[1][0] = 1128ns;
slave_timing[0][160+11].t_rxd1[0][2] = 794ns;
slave_timing[0][160+11].t_rxd1[2][0] = 1412ns;
slave_timing[0][160+11].t_rxd2[0][2] = 1326ns;
slave_timing[0][160+11].t_rxd2[2][0] = 834ns;
slave_timing[0][160+11].t_rxd2[1][2] = 1036ns;
slave_timing[0][160+11].t_rxd2[2][1] = 1141ns;

slave_timing[0][160+12].info_corner          = 2;
slave_timing[0][160+12].info_temp__j__       = -40;
slave_timing[0][160+12].info_i__quite_rec__  = 0.003000000;
slave_timing[0][160+12].info_dtr__ib__       = -1;
slave_timing[0][160+12].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+12].info_i__max_slave__  = 0.023000000;
slave_timing[0][160+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][160+12].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+12].t_rxd1[0][1] = 1164ns;
slave_timing[0][160+12].t_rxd1[1][0] = 1188ns;
slave_timing[0][160+12].t_rxd1[0][2] = 860ns;
slave_timing[0][160+12].t_rxd1[2][0] = 1468ns;
slave_timing[0][160+12].t_rxd2[0][2] = 1380ns;
slave_timing[0][160+12].t_rxd2[2][0] = 839ns;
slave_timing[0][160+12].t_rxd2[1][2] = 1082ns;
slave_timing[0][160+12].t_rxd2[2][1] = 1119ns;

slave_timing[0][160+13].info_corner          = 2;
slave_timing[0][160+13].info_temp__j__       = -40;
slave_timing[0][160+13].info_i__quite_rec__  = 0.003000000;
slave_timing[0][160+13].info_dtr__ib__       = -1;
slave_timing[0][160+13].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+13].info_i__max_slave__  = 0.025000000;
slave_timing[0][160+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][160+13].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+13].t_rxd1[0][1] = 1112ns;
slave_timing[0][160+13].t_rxd1[1][0] = 1219ns;
slave_timing[0][160+13].t_rxd1[0][2] = 835ns;
slave_timing[0][160+13].t_rxd1[2][0] = 1498ns;
slave_timing[0][160+13].t_rxd2[0][2] = 1282ns;
slave_timing[0][160+13].t_rxd2[2][0] = 891ns;
slave_timing[0][160+13].t_rxd2[1][2] = 960ns;
slave_timing[0][160+13].t_rxd2[2][1] = 1250ns;

slave_timing[0][160+14].info_corner          = 2;
slave_timing[0][160+14].info_temp__j__       = -40;
slave_timing[0][160+14].info_i__quite_rec__  = 0.003000000;
slave_timing[0][160+14].info_dtr__ib__       = 1;
slave_timing[0][160+14].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+14].info_i__max_slave__  = 0.023000000;
slave_timing[0][160+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][160+14].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+14].t_rxd1[0][1] = 1195ns;
slave_timing[0][160+14].t_rxd1[1][0] = 1154ns;
slave_timing[0][160+14].t_rxd1[0][2] = 871ns;
slave_timing[0][160+14].t_rxd1[2][0] = 1437ns;
slave_timing[0][160+14].t_rxd2[0][2] = 1471ns;
slave_timing[0][160+14].t_rxd2[2][0] = 790ns;
slave_timing[0][160+14].t_rxd2[1][2] = 1187ns;
slave_timing[0][160+14].t_rxd2[2][1] = 1027ns;

slave_timing[0][160+15].info_corner          = 2;
slave_timing[0][160+15].info_temp__j__       = -40;
slave_timing[0][160+15].info_i__quite_rec__  = 0.003000000;
slave_timing[0][160+15].info_dtr__ib__       = 1;
slave_timing[0][160+15].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+15].info_i__max_slave__  = 0.025000000;
slave_timing[0][160+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][160+15].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+15].t_rxd1[0][1] = 1140ns;
slave_timing[0][160+15].t_rxd1[1][0] = 1192ns;
slave_timing[0][160+15].t_rxd1[0][2] = 843ns;
slave_timing[0][160+15].t_rxd1[2][0] = 1468ns;
slave_timing[0][160+15].t_rxd2[0][2] = 1346ns;
slave_timing[0][160+15].t_rxd2[2][0] = 849ns;
slave_timing[0][160+15].t_rxd2[1][2] = 1043ns;
slave_timing[0][160+15].t_rxd2[2][1] = 1151ns;

slave_timing[0][160+16].info_corner          = 2;
slave_timing[0][160+16].info_temp__j__       = -40;
slave_timing[0][160+16].info_i__quite_rec__  = 0.000000000;
slave_timing[0][160+16].info_dtr__ib__       = -1;
slave_timing[0][160+16].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+16].info_i__max_slave__  = 0.023000000;
slave_timing[0][160+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][160+16].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+16].t_rxd1[0][1] = 1101ns;
slave_timing[0][160+16].t_rxd1[1][0] = 1113ns;
slave_timing[0][160+16].t_rxd1[0][2] = 808ns;
slave_timing[0][160+16].t_rxd1[2][0] = 1398ns;
slave_timing[0][160+16].t_rxd2[0][2] = 1364ns;
slave_timing[0][160+16].t_rxd2[2][0] = 814ns;
slave_timing[0][160+16].t_rxd2[1][2] = 1081ns;
slave_timing[0][160+16].t_rxd2[2][1] = 1099ns;

slave_timing[0][160+17].info_corner          = 2;
slave_timing[0][160+17].info_temp__j__       = -40;
slave_timing[0][160+17].info_i__quite_rec__  = 0.000000000;
slave_timing[0][160+17].info_dtr__ib__       = -1;
slave_timing[0][160+17].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+17].info_i__max_slave__  = 0.025000000;
slave_timing[0][160+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][160+17].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+17].t_rxd1[0][1] = 1051ns;
slave_timing[0][160+17].t_rxd1[1][0] = 1145ns;
slave_timing[0][160+17].t_rxd1[0][2] = 785ns;
slave_timing[0][160+17].t_rxd1[2][0] = 1429ns;
slave_timing[0][160+17].t_rxd2[0][2] = 1264ns;
slave_timing[0][160+17].t_rxd2[2][0] = 869ns;
slave_timing[0][160+17].t_rxd2[1][2] = 952ns;
slave_timing[0][160+17].t_rxd2[2][1] = 1233ns;

slave_timing[0][160+18].info_corner          = 2;
slave_timing[0][160+18].info_temp__j__       = -40;
slave_timing[0][160+18].info_i__quite_rec__  = 0.000000000;
slave_timing[0][160+18].info_dtr__ib__       = 1;
slave_timing[0][160+18].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+18].info_i__max_slave__  = 0.023000000;
slave_timing[0][160+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][160+18].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+18].t_rxd1[0][1] = 1140ns;
slave_timing[0][160+18].t_rxd1[1][0] = 1080ns;
slave_timing[0][160+18].t_rxd1[0][2] = 827ns;
slave_timing[0][160+18].t_rxd1[2][0] = 1371ns;
slave_timing[0][160+18].t_rxd2[0][2] = 1464ns;
slave_timing[0][160+18].t_rxd2[2][0] = 764ns;
slave_timing[0][160+18].t_rxd2[1][2] = 1191ns;
slave_timing[0][160+18].t_rxd2[2][1] = 998ns;

slave_timing[0][160+19].info_corner          = 2;
slave_timing[0][160+19].info_temp__j__       = -40;
slave_timing[0][160+19].info_i__quite_rec__  = 0.000000000;
slave_timing[0][160+19].info_dtr__ib__       = 1;
slave_timing[0][160+19].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+19].info_i__max_slave__  = 0.025000000;
slave_timing[0][160+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][160+19].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+19].t_rxd1[0][1] = 1086ns;
slave_timing[0][160+19].t_rxd1[1][0] = 1118ns;
slave_timing[0][160+19].t_rxd1[0][2] = 802ns;
slave_timing[0][160+19].t_rxd1[2][0] = 1403ns;
slave_timing[0][160+19].t_rxd2[0][2] = 1336ns;
slave_timing[0][160+19].t_rxd2[2][0] = 825ns;
slave_timing[0][160+19].t_rxd2[1][2] = 1046ns;
slave_timing[0][160+19].t_rxd2[2][1] = 1125ns;

slave_timing[0][160+20].info_corner          = 2;
slave_timing[0][160+20].info_temp__j__       = -40;
slave_timing[0][160+20].info_i__quite_rec__  = 0.000000000;
slave_timing[0][160+20].info_dtr__ib__       = -1;
slave_timing[0][160+20].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+20].info_i__max_slave__  = 0.023000000;
slave_timing[0][160+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][160+20].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+20].t_rxd1[0][1] = 1179ns;
slave_timing[0][160+20].t_rxd1[1][0] = 1181ns;
slave_timing[0][160+20].t_rxd1[0][2] = 868ns;
slave_timing[0][160+20].t_rxd1[2][0] = 1463ns;
slave_timing[0][160+20].t_rxd2[0][2] = 1389ns;
slave_timing[0][160+20].t_rxd2[2][0] = 832ns;
slave_timing[0][160+20].t_rxd2[1][2] = 1090ns;
slave_timing[0][160+20].t_rxd2[2][1] = 1108ns;

slave_timing[0][160+21].info_corner          = 2;
slave_timing[0][160+21].info_temp__j__       = -40;
slave_timing[0][160+21].info_i__quite_rec__  = 0.000000000;
slave_timing[0][160+21].info_dtr__ib__       = -1;
slave_timing[0][160+21].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+21].info_i__max_slave__  = 0.025000000;
slave_timing[0][160+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][160+21].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+21].t_rxd1[0][1] = 1126ns;
slave_timing[0][160+21].t_rxd1[1][0] = 1217ns;
slave_timing[0][160+21].t_rxd1[0][2] = 844ns;
slave_timing[0][160+21].t_rxd1[2][0] = 1492ns;
slave_timing[0][160+21].t_rxd2[0][2] = 1289ns;
slave_timing[0][160+21].t_rxd2[2][0] = 885ns;
slave_timing[0][160+21].t_rxd2[1][2] = 966ns;
slave_timing[0][160+21].t_rxd2[2][1] = 1240ns;

slave_timing[0][160+22].info_corner          = 2;
slave_timing[0][160+22].info_temp__j__       = -40;
slave_timing[0][160+22].info_i__quite_rec__  = 0.000000000;
slave_timing[0][160+22].info_dtr__ib__       = 1;
slave_timing[0][160+22].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+22].info_i__max_slave__  = 0.023000000;
slave_timing[0][160+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][160+22].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+22].t_rxd1[0][1] = 1213ns;
slave_timing[0][160+22].t_rxd1[1][0] = 1146ns;
slave_timing[0][160+22].t_rxd1[0][2] = 880ns;
slave_timing[0][160+22].t_rxd1[2][0] = 1433ns;
slave_timing[0][160+22].t_rxd2[0][2] = 1483ns;
slave_timing[0][160+22].t_rxd2[2][0] = 782ns;
slave_timing[0][160+22].t_rxd2[1][2] = 1200ns;
slave_timing[0][160+22].t_rxd2[2][1] = 1010ns;

slave_timing[0][160+23].info_corner          = 2;
slave_timing[0][160+23].info_temp__j__       = -40;
slave_timing[0][160+23].info_i__quite_rec__  = 0.000000000;
slave_timing[0][160+23].info_dtr__ib__       = 1;
slave_timing[0][160+23].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+23].info_i__max_slave__  = 0.025000000;
slave_timing[0][160+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][160+23].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+23].t_rxd1[0][1] = 1155ns;
slave_timing[0][160+23].t_rxd1[1][0] = 1183ns;
slave_timing[0][160+23].t_rxd1[0][2] = 856ns;
slave_timing[0][160+23].t_rxd1[2][0] = 1463ns;
slave_timing[0][160+23].t_rxd2[0][2] = 1356ns;
slave_timing[0][160+23].t_rxd2[2][0] = 842ns;
slave_timing[0][160+23].t_rxd2[1][2] = 1056ns;
slave_timing[0][160+23].t_rxd2[2][1] = 1133ns;

slave_timing[0][160+24].info_corner          = 2;
slave_timing[0][160+24].info_temp__j__       = -40;
slave_timing[0][160+24].info_i__quite_rec__  = 0.040000000;
slave_timing[0][160+24].info_dtr__ib__       = -1;
slave_timing[0][160+24].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+24].info_i__max_slave__  = 0.023000000;
slave_timing[0][160+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][160+24].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+24].t_rxd1[0][1] = 1093ns;
slave_timing[0][160+24].t_rxd1[1][0] = 1103ns;
slave_timing[0][160+24].t_rxd1[0][2] = 805ns;
slave_timing[0][160+24].t_rxd1[2][0] = 1389ns;
slave_timing[0][160+24].t_rxd2[0][2] = 1363ns;
slave_timing[0][160+24].t_rxd2[2][0] = 813ns;
slave_timing[0][160+24].t_rxd2[1][2] = 1080ns;
slave_timing[0][160+24].t_rxd2[2][1] = 1097ns;

slave_timing[0][160+25].info_corner          = 2;
slave_timing[0][160+25].info_temp__j__       = -40;
slave_timing[0][160+25].info_i__quite_rec__  = 0.040000000;
slave_timing[0][160+25].info_dtr__ib__       = -1;
slave_timing[0][160+25].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+25].info_i__max_slave__  = 0.025000000;
slave_timing[0][160+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][160+25].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+25].t_rxd1[0][1] = 1046ns;
slave_timing[0][160+25].t_rxd1[1][0] = 1139ns;
slave_timing[0][160+25].t_rxd1[0][2] = 781ns;
slave_timing[0][160+25].t_rxd1[2][0] = 1419ns;
slave_timing[0][160+25].t_rxd2[0][2] = 1262ns;
slave_timing[0][160+25].t_rxd2[2][0] = 867ns;
slave_timing[0][160+25].t_rxd2[1][2] = 956ns;
slave_timing[0][160+25].t_rxd2[2][1] = 1229ns;

slave_timing[0][160+26].info_corner          = 2;
slave_timing[0][160+26].info_temp__j__       = -40;
slave_timing[0][160+26].info_i__quite_rec__  = 0.040000000;
slave_timing[0][160+26].info_dtr__ib__       = 1;
slave_timing[0][160+26].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+26].info_i__max_slave__  = 0.023000000;
slave_timing[0][160+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][160+26].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+26].t_rxd1[0][1] = 1125ns;
slave_timing[0][160+26].t_rxd1[1][0] = 1080ns;
slave_timing[0][160+26].t_rxd1[0][2] = 819ns;
slave_timing[0][160+26].t_rxd1[2][0] = 1371ns;
slave_timing[0][160+26].t_rxd2[0][2] = 1455ns;
slave_timing[0][160+26].t_rxd2[2][0] = 769ns;
slave_timing[0][160+26].t_rxd2[1][2] = 1185ns;
slave_timing[0][160+26].t_rxd2[2][1] = 1007ns;

slave_timing[0][160+27].info_corner          = 2;
slave_timing[0][160+27].info_temp__j__       = -40;
slave_timing[0][160+27].info_i__quite_rec__  = 0.040000000;
slave_timing[0][160+27].info_dtr__ib__       = 1;
slave_timing[0][160+27].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+27].info_i__max_slave__  = 0.025000000;
slave_timing[0][160+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][160+27].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+27].t_rxd1[0][1] = 1070ns;
slave_timing[0][160+27].t_rxd1[1][0] = 1116ns;
slave_timing[0][160+27].t_rxd1[0][2] = 793ns;
slave_timing[0][160+27].t_rxd1[2][0] = 1403ns;
slave_timing[0][160+27].t_rxd2[0][2] = 1328ns;
slave_timing[0][160+27].t_rxd2[2][0] = 828ns;
slave_timing[0][160+27].t_rxd2[1][2] = 1042ns;
slave_timing[0][160+27].t_rxd2[2][1] = 1132ns;

slave_timing[0][160+28].info_corner          = 2;
slave_timing[0][160+28].info_temp__j__       = -40;
slave_timing[0][160+28].info_i__quite_rec__  = 0.040000000;
slave_timing[0][160+28].info_dtr__ib__       = -1;
slave_timing[0][160+28].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+28].info_i__max_slave__  = 0.023000000;
slave_timing[0][160+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][160+28].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+28].t_rxd1[0][1] = 1132ns;
slave_timing[0][160+28].t_rxd1[1][0] = 1144ns;
slave_timing[0][160+28].t_rxd1[0][2] = 841ns;
slave_timing[0][160+28].t_rxd1[2][0] = 1423ns;
slave_timing[0][160+28].t_rxd2[0][2] = 1377ns;
slave_timing[0][160+28].t_rxd2[2][0] = 832ns;
slave_timing[0][160+28].t_rxd2[1][2] = 1093ns;
slave_timing[0][160+28].t_rxd2[2][1] = 1106ns;

slave_timing[0][160+29].info_corner          = 2;
slave_timing[0][160+29].info_temp__j__       = -40;
slave_timing[0][160+29].info_i__quite_rec__  = 0.040000000;
slave_timing[0][160+29].info_dtr__ib__       = -1;
slave_timing[0][160+29].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+29].info_i__max_slave__  = 0.025000000;
slave_timing[0][160+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][160+29].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+29].t_rxd1[0][1] = 1085ns;
slave_timing[0][160+29].t_rxd1[1][0] = 1178ns;
slave_timing[0][160+29].t_rxd1[0][2] = 815ns;
slave_timing[0][160+29].t_rxd1[2][0] = 1453ns;
slave_timing[0][160+29].t_rxd2[0][2] = 1277ns;
slave_timing[0][160+29].t_rxd2[2][0] = 885ns;
slave_timing[0][160+29].t_rxd2[1][2] = 968ns;
slave_timing[0][160+29].t_rxd2[2][1] = 1236ns;

slave_timing[0][160+30].info_corner          = 2;
slave_timing[0][160+30].info_temp__j__       = -40;
slave_timing[0][160+30].info_i__quite_rec__  = 0.040000000;
slave_timing[0][160+30].info_dtr__ib__       = 1;
slave_timing[0][160+30].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+30].info_i__max_slave__  = 0.023000000;
slave_timing[0][160+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][160+30].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+30].t_rxd1[0][1] = 1160ns;
slave_timing[0][160+30].t_rxd1[1][0] = 1117ns;
slave_timing[0][160+30].t_rxd1[0][2] = 850ns;
slave_timing[0][160+30].t_rxd1[2][0] = 1402ns;
slave_timing[0][160+30].t_rxd2[0][2] = 1463ns;
slave_timing[0][160+30].t_rxd2[2][0] = 784ns;
slave_timing[0][160+30].t_rxd2[1][2] = 1194ns;
slave_timing[0][160+30].t_rxd2[2][1] = 1016ns;

slave_timing[0][160+31].info_corner          = 2;
slave_timing[0][160+31].info_temp__j__       = -40;
slave_timing[0][160+31].info_i__quite_rec__  = 0.040000000;
slave_timing[0][160+31].info_dtr__ib__       = 1;
slave_timing[0][160+31].info_i__offset_rec__ = 0.000000000;
slave_timing[0][160+31].info_i__max_slave__  = 0.025000000;
slave_timing[0][160+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][160+31].info_r__dsi_bus__    = 5.000;

slave_timing[0][160+31].t_rxd1[0][1] = 1110ns;
slave_timing[0][160+31].t_rxd1[1][0] = 1156ns;
slave_timing[0][160+31].t_rxd1[0][2] = 828ns;
slave_timing[0][160+31].t_rxd1[2][0] = 1433ns;
slave_timing[0][160+31].t_rxd2[0][2] = 1341ns;
slave_timing[0][160+31].t_rxd2[2][0] = 843ns;
slave_timing[0][160+31].t_rxd2[1][2] = 1052ns;
slave_timing[0][160+31].t_rxd2[2][1] = 1140ns;


/*==================================================
 *  Copyright (c) 2023 Elmos SE
 *  Author: stove
 *  Description : Note: This file has been generated automatically by stove
 *                Note: This file should not be modified manually.
 *                test interface definition for TEST_WS
 *==================================================*/
interface tmr_ws_if;



modport master (
);

modport slave (
);

modport iomux (
);



endinterface

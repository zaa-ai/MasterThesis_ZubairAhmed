virtual clk_reset_if vif_clk_rst;

buffer_writer_action_e action;

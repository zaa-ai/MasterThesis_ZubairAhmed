
slave_timing[0][192+0].info_corner          = 3;
slave_timing[0][192+0].info_temp__j__       = -40;
slave_timing[0][192+0].info_i__quite_rec__  = 0.006000000;
slave_timing[0][192+0].info_dtr__ib__       = -1;
slave_timing[0][192+0].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+0].info_i__max_slave__  = 0.023000000;
slave_timing[0][192+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][192+0].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+0].t_rxd1[0][1] = 1096ns;
slave_timing[0][192+0].t_rxd1[1][0] = 1120ns;
slave_timing[0][192+0].t_rxd1[0][2] = 809ns;
slave_timing[0][192+0].t_rxd1[2][0] = 1408ns;
slave_timing[0][192+0].t_rxd2[0][2] = 1361ns;
slave_timing[0][192+0].t_rxd2[2][0] = 821ns;
slave_timing[0][192+0].t_rxd2[1][2] = 1068ns;
slave_timing[0][192+0].t_rxd2[2][1] = 1112ns;

slave_timing[0][192+1].info_corner          = 3;
slave_timing[0][192+1].info_temp__j__       = -40;
slave_timing[0][192+1].info_i__quite_rec__  = 0.006000000;
slave_timing[0][192+1].info_dtr__ib__       = -1;
slave_timing[0][192+1].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+1].info_i__max_slave__  = 0.025000000;
slave_timing[0][192+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][192+1].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+1].t_rxd1[0][1] = 1048ns;
slave_timing[0][192+1].t_rxd1[1][0] = 1155ns;
slave_timing[0][192+1].t_rxd1[0][2] = 783ns;
slave_timing[0][192+1].t_rxd1[2][0] = 1439ns;
slave_timing[0][192+1].t_rxd2[0][2] = 1262ns;
slave_timing[0][192+1].t_rxd2[2][0] = 875ns;
slave_timing[0][192+1].t_rxd2[1][2] = 942ns;
slave_timing[0][192+1].t_rxd2[2][1] = 1251ns;

slave_timing[0][192+2].info_corner          = 3;
slave_timing[0][192+2].info_temp__j__       = -40;
slave_timing[0][192+2].info_i__quite_rec__  = 0.006000000;
slave_timing[0][192+2].info_dtr__ib__       = 1;
slave_timing[0][192+2].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+2].info_i__max_slave__  = 0.023000000;
slave_timing[0][192+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][192+2].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+2].t_rxd1[0][1] = 1130ns;
slave_timing[0][192+2].t_rxd1[1][0] = 1088ns;
slave_timing[0][192+2].t_rxd1[0][2] = 825ns;
slave_timing[0][192+2].t_rxd1[2][0] = 1384ns;
slave_timing[0][192+2].t_rxd2[0][2] = 1455ns;
slave_timing[0][192+2].t_rxd2[2][0] = 775ns;
slave_timing[0][192+2].t_rxd2[1][2] = 1176ns;
slave_timing[0][192+2].t_rxd2[2][1] = 1020ns;

slave_timing[0][192+3].info_corner          = 3;
slave_timing[0][192+3].info_temp__j__       = -40;
slave_timing[0][192+3].info_i__quite_rec__  = 0.006000000;
slave_timing[0][192+3].info_dtr__ib__       = 1;
slave_timing[0][192+3].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+3].info_i__max_slave__  = 0.025000000;
slave_timing[0][192+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][192+3].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+3].t_rxd1[0][1] = 1077ns;
slave_timing[0][192+3].t_rxd1[1][0] = 1128ns;
slave_timing[0][192+3].t_rxd1[0][2] = 799ns;
slave_timing[0][192+3].t_rxd1[2][0] = 1416ns;
slave_timing[0][192+3].t_rxd2[0][2] = 1329ns;
slave_timing[0][192+3].t_rxd2[2][0] = 835ns;
slave_timing[0][192+3].t_rxd2[1][2] = 1032ns;
slave_timing[0][192+3].t_rxd2[2][1] = 1145ns;

slave_timing[0][192+4].info_corner          = 3;
slave_timing[0][192+4].info_temp__j__       = -40;
slave_timing[0][192+4].info_i__quite_rec__  = 0.006000000;
slave_timing[0][192+4].info_dtr__ib__       = -1;
slave_timing[0][192+4].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+4].info_i__max_slave__  = 0.023000000;
slave_timing[0][192+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][192+4].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+4].t_rxd1[0][1] = 1180ns;
slave_timing[0][192+4].t_rxd1[1][0] = 1197ns;
slave_timing[0][192+4].t_rxd1[0][2] = 871ns;
slave_timing[0][192+4].t_rxd1[2][0] = 1481ns;
slave_timing[0][192+4].t_rxd2[0][2] = 1390ns;
slave_timing[0][192+4].t_rxd2[2][0] = 843ns;
slave_timing[0][192+4].t_rxd2[1][2] = 1082ns;
slave_timing[0][192+4].t_rxd2[2][1] = 1129ns;

slave_timing[0][192+5].info_corner          = 3;
slave_timing[0][192+5].info_temp__j__       = -40;
slave_timing[0][192+5].info_i__quite_rec__  = 0.006000000;
slave_timing[0][192+5].info_dtr__ib__       = -1;
slave_timing[0][192+5].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+5].info_i__max_slave__  = 0.025000000;
slave_timing[0][192+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][192+5].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+5].t_rxd1[0][1] = 1128ns;
slave_timing[0][192+5].t_rxd1[1][0] = 1233ns;
slave_timing[0][192+5].t_rxd1[0][2] = 845ns;
slave_timing[0][192+5].t_rxd1[2][0] = 1510ns;
slave_timing[0][192+5].t_rxd2[0][2] = 1292ns;
slave_timing[0][192+5].t_rxd2[2][0] = 897ns;
slave_timing[0][192+5].t_rxd2[1][2] = 961ns;
slave_timing[0][192+5].t_rxd2[2][1] = 1264ns;

slave_timing[0][192+6].info_corner          = 3;
slave_timing[0][192+6].info_temp__j__       = -40;
slave_timing[0][192+6].info_i__quite_rec__  = 0.006000000;
slave_timing[0][192+6].info_dtr__ib__       = 1;
slave_timing[0][192+6].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+6].info_i__max_slave__  = 0.023000000;
slave_timing[0][192+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][192+6].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+6].t_rxd1[0][1] = 1208ns;
slave_timing[0][192+6].t_rxd1[1][0] = 1161ns;
slave_timing[0][192+6].t_rxd1[0][2] = 882ns;
slave_timing[0][192+6].t_rxd1[2][0] = 1450ns;
slave_timing[0][192+6].t_rxd2[0][2] = 1480ns;
slave_timing[0][192+6].t_rxd2[2][0] = 795ns;
slave_timing[0][192+6].t_rxd2[1][2] = 1188ns;
slave_timing[0][192+6].t_rxd2[2][1] = 1034ns;

slave_timing[0][192+7].info_corner          = 3;
slave_timing[0][192+7].info_temp__j__       = -40;
slave_timing[0][192+7].info_i__quite_rec__  = 0.006000000;
slave_timing[0][192+7].info_dtr__ib__       = 1;
slave_timing[0][192+7].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+7].info_i__max_slave__  = 0.025000000;
slave_timing[0][192+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][192+7].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+7].t_rxd1[0][1] = 1154ns;
slave_timing[0][192+7].t_rxd1[1][0] = 1199ns;
slave_timing[0][192+7].t_rxd1[0][2] = 855ns;
slave_timing[0][192+7].t_rxd1[2][0] = 1480ns;
slave_timing[0][192+7].t_rxd2[0][2] = 1354ns;
slave_timing[0][192+7].t_rxd2[2][0] = 853ns;
slave_timing[0][192+7].t_rxd2[1][2] = 1047ns;
slave_timing[0][192+7].t_rxd2[2][1] = 1158ns;

slave_timing[0][192+8].info_corner          = 3;
slave_timing[0][192+8].info_temp__j__       = -40;
slave_timing[0][192+8].info_i__quite_rec__  = 0.003000000;
slave_timing[0][192+8].info_dtr__ib__       = -1;
slave_timing[0][192+8].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+8].info_i__max_slave__  = 0.023000000;
slave_timing[0][192+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][192+8].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+8].t_rxd1[0][1] = 1089ns;
slave_timing[0][192+8].t_rxd1[1][0] = 1124ns;
slave_timing[0][192+8].t_rxd1[0][2] = 806ns;
slave_timing[0][192+8].t_rxd1[2][0] = 1418ns;
slave_timing[0][192+8].t_rxd2[0][2] = 1355ns;
slave_timing[0][192+8].t_rxd2[2][0] = 823ns;
slave_timing[0][192+8].t_rxd2[1][2] = 1061ns;
slave_timing[0][192+8].t_rxd2[2][1] = 1116ns;

slave_timing[0][192+9].info_corner          = 3;
slave_timing[0][192+9].info_temp__j__       = -40;
slave_timing[0][192+9].info_i__quite_rec__  = 0.003000000;
slave_timing[0][192+9].info_dtr__ib__       = -1;
slave_timing[0][192+9].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+9].info_i__max_slave__  = 0.025000000;
slave_timing[0][192+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][192+9].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+9].t_rxd1[0][1] = 1044ns;
slave_timing[0][192+9].t_rxd1[1][0] = 1163ns;
slave_timing[0][192+9].t_rxd1[0][2] = 782ns;
slave_timing[0][192+9].t_rxd1[2][0] = 1448ns;
slave_timing[0][192+9].t_rxd2[0][2] = 1258ns;
slave_timing[0][192+9].t_rxd2[2][0] = 875ns;
slave_timing[0][192+9].t_rxd2[1][2] = 937ns;
slave_timing[0][192+9].t_rxd2[2][1] = 1255ns;

slave_timing[0][192+10].info_corner          = 3;
slave_timing[0][192+10].info_temp__j__       = -40;
slave_timing[0][192+10].info_i__quite_rec__  = 0.003000000;
slave_timing[0][192+10].info_dtr__ib__       = 1;
slave_timing[0][192+10].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+10].info_i__max_slave__  = 0.023000000;
slave_timing[0][192+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][192+10].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+10].t_rxd1[0][1] = 1125ns;
slave_timing[0][192+10].t_rxd1[1][0] = 1095ns;
slave_timing[0][192+10].t_rxd1[0][2] = 810ns;
slave_timing[0][192+10].t_rxd1[2][0] = 1388ns;
slave_timing[0][192+10].t_rxd2[0][2] = 1429ns;
slave_timing[0][192+10].t_rxd2[2][0] = 779ns;
slave_timing[0][192+10].t_rxd2[1][2] = 1171ns;
slave_timing[0][192+10].t_rxd2[2][1] = 1022ns;

slave_timing[0][192+11].info_corner          = 3;
slave_timing[0][192+11].info_temp__j__       = -40;
slave_timing[0][192+11].info_i__quite_rec__  = 0.003000000;
slave_timing[0][192+11].info_dtr__ib__       = 1;
slave_timing[0][192+11].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+11].info_i__max_slave__  = 0.025000000;
slave_timing[0][192+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][192+11].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+11].t_rxd1[0][1] = 1074ns;
slave_timing[0][192+11].t_rxd1[1][0] = 1129ns;
slave_timing[0][192+11].t_rxd1[0][2] = 798ns;
slave_timing[0][192+11].t_rxd1[2][0] = 1419ns;
slave_timing[0][192+11].t_rxd2[0][2] = 1328ns;
slave_timing[0][192+11].t_rxd2[2][0] = 837ns;
slave_timing[0][192+11].t_rxd2[1][2] = 1028ns;
slave_timing[0][192+11].t_rxd2[2][1] = 1148ns;

slave_timing[0][192+12].info_corner          = 3;
slave_timing[0][192+12].info_temp__j__       = -40;
slave_timing[0][192+12].info_i__quite_rec__  = 0.003000000;
slave_timing[0][192+12].info_dtr__ib__       = -1;
slave_timing[0][192+12].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+12].info_i__max_slave__  = 0.023000000;
slave_timing[0][192+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][192+12].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+12].t_rxd1[0][1] = 1178ns;
slave_timing[0][192+12].t_rxd1[1][0] = 1207ns;
slave_timing[0][192+12].t_rxd1[0][2] = 871ns;
slave_timing[0][192+12].t_rxd1[2][0] = 1490ns;
slave_timing[0][192+12].t_rxd2[0][2] = 1383ns;
slave_timing[0][192+12].t_rxd2[2][0] = 843ns;
slave_timing[0][192+12].t_rxd2[1][2] = 1092ns;
slave_timing[0][192+12].t_rxd2[2][1] = 1112ns;

slave_timing[0][192+13].info_corner          = 3;
slave_timing[0][192+13].info_temp__j__       = -40;
slave_timing[0][192+13].info_i__quite_rec__  = 0.003000000;
slave_timing[0][192+13].info_dtr__ib__       = -1;
slave_timing[0][192+13].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+13].info_i__max_slave__  = 0.025000000;
slave_timing[0][192+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][192+13].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+13].t_rxd1[0][1] = 1129ns;
slave_timing[0][192+13].t_rxd1[1][0] = 1244ns;
slave_timing[0][192+13].t_rxd1[0][2] = 849ns;
slave_timing[0][192+13].t_rxd1[2][0] = 1521ns;
slave_timing[0][192+13].t_rxd2[0][2] = 1290ns;
slave_timing[0][192+13].t_rxd2[2][0] = 897ns;
slave_timing[0][192+13].t_rxd2[1][2] = 953ns;
slave_timing[0][192+13].t_rxd2[2][1] = 1264ns;

slave_timing[0][192+14].info_corner          = 3;
slave_timing[0][192+14].info_temp__j__       = -40;
slave_timing[0][192+14].info_i__quite_rec__  = 0.003000000;
slave_timing[0][192+14].info_dtr__ib__       = 1;
slave_timing[0][192+14].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+14].info_i__max_slave__  = 0.023000000;
slave_timing[0][192+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][192+14].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+14].t_rxd1[0][1] = 1206ns;
slave_timing[0][192+14].t_rxd1[1][0] = 1163ns;
slave_timing[0][192+14].t_rxd1[0][2] = 881ns;
slave_timing[0][192+14].t_rxd1[2][0] = 1454ns;
slave_timing[0][192+14].t_rxd2[0][2] = 1475ns;
slave_timing[0][192+14].t_rxd2[2][0] = 794ns;
slave_timing[0][192+14].t_rxd2[1][2] = 1182ns;
slave_timing[0][192+14].t_rxd2[2][1] = 1036ns;

slave_timing[0][192+15].info_corner          = 3;
slave_timing[0][192+15].info_temp__j__       = -40;
slave_timing[0][192+15].info_i__quite_rec__  = 0.003000000;
slave_timing[0][192+15].info_dtr__ib__       = 1;
slave_timing[0][192+15].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+15].info_i__max_slave__  = 0.025000000;
slave_timing[0][192+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][192+15].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+15].t_rxd1[0][1] = 1151ns;
slave_timing[0][192+15].t_rxd1[1][0] = 1204ns;
slave_timing[0][192+15].t_rxd1[0][2] = 847ns;
slave_timing[0][192+15].t_rxd1[2][0] = 1485ns;
slave_timing[0][192+15].t_rxd2[0][2] = 1339ns;
slave_timing[0][192+15].t_rxd2[2][0] = 855ns;
slave_timing[0][192+15].t_rxd2[1][2] = 1041ns;
slave_timing[0][192+15].t_rxd2[2][1] = 1161ns;

slave_timing[0][192+16].info_corner          = 3;
slave_timing[0][192+16].info_temp__j__       = -40;
slave_timing[0][192+16].info_i__quite_rec__  = 0.000000000;
slave_timing[0][192+16].info_dtr__ib__       = -1;
slave_timing[0][192+16].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+16].info_i__max_slave__  = 0.023000000;
slave_timing[0][192+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][192+16].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+16].t_rxd1[0][1] = 1104ns;
slave_timing[0][192+16].t_rxd1[1][0] = 1112ns;
slave_timing[0][192+16].t_rxd1[0][2] = 812ns;
slave_timing[0][192+16].t_rxd1[2][0] = 1403ns;
slave_timing[0][192+16].t_rxd2[0][2] = 1365ns;
slave_timing[0][192+16].t_rxd2[2][0] = 814ns;
slave_timing[0][192+16].t_rxd2[1][2] = 1075ns;
slave_timing[0][192+16].t_rxd2[2][1] = 1106ns;

slave_timing[0][192+17].info_corner          = 3;
slave_timing[0][192+17].info_temp__j__       = -40;
slave_timing[0][192+17].info_i__quite_rec__  = 0.000000000;
slave_timing[0][192+17].info_dtr__ib__       = -1;
slave_timing[0][192+17].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+17].info_i__max_slave__  = 0.025000000;
slave_timing[0][192+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][192+17].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+17].t_rxd1[0][1] = 1056ns;
slave_timing[0][192+17].t_rxd1[1][0] = 1151ns;
slave_timing[0][192+17].t_rxd1[0][2] = 787ns;
slave_timing[0][192+17].t_rxd1[2][0] = 1436ns;
slave_timing[0][192+17].t_rxd2[0][2] = 1266ns;
slave_timing[0][192+17].t_rxd2[2][0] = 872ns;
slave_timing[0][192+17].t_rxd2[1][2] = 952ns;
slave_timing[0][192+17].t_rxd2[2][1] = 1244ns;

slave_timing[0][192+18].info_corner          = 3;
slave_timing[0][192+18].info_temp__j__       = -40;
slave_timing[0][192+18].info_i__quite_rec__  = 0.000000000;
slave_timing[0][192+18].info_dtr__ib__       = 1;
slave_timing[0][192+18].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+18].info_i__max_slave__  = 0.023000000;
slave_timing[0][192+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][192+18].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+18].t_rxd1[0][1] = 1142ns;
slave_timing[0][192+18].t_rxd1[1][0] = 1083ns;
slave_timing[0][192+18].t_rxd1[0][2] = 829ns;
slave_timing[0][192+18].t_rxd1[2][0] = 1375ns;
slave_timing[0][192+18].t_rxd2[0][2] = 1462ns;
slave_timing[0][192+18].t_rxd2[2][0] = 767ns;
slave_timing[0][192+18].t_rxd2[1][2] = 1188ns;
slave_timing[0][192+18].t_rxd2[2][1] = 1009ns;

slave_timing[0][192+19].info_corner          = 3;
slave_timing[0][192+19].info_temp__j__       = -40;
slave_timing[0][192+19].info_i__quite_rec__  = 0.000000000;
slave_timing[0][192+19].info_dtr__ib__       = 1;
slave_timing[0][192+19].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+19].info_i__max_slave__  = 0.025000000;
slave_timing[0][192+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][192+19].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+19].t_rxd1[0][1] = 1088ns;
slave_timing[0][192+19].t_rxd1[1][0] = 1120ns;
slave_timing[0][192+19].t_rxd1[0][2] = 805ns;
slave_timing[0][192+19].t_rxd1[2][0] = 1409ns;
slave_timing[0][192+19].t_rxd2[0][2] = 1337ns;
slave_timing[0][192+19].t_rxd2[2][0] = 829ns;
slave_timing[0][192+19].t_rxd2[1][2] = 1039ns;
slave_timing[0][192+19].t_rxd2[2][1] = 1136ns;

slave_timing[0][192+20].info_corner          = 3;
slave_timing[0][192+20].info_temp__j__       = -40;
slave_timing[0][192+20].info_i__quite_rec__  = 0.000000000;
slave_timing[0][192+20].info_dtr__ib__       = -1;
slave_timing[0][192+20].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+20].info_i__max_slave__  = 0.023000000;
slave_timing[0][192+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][192+20].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+20].t_rxd1[0][1] = 1197ns;
slave_timing[0][192+20].t_rxd1[1][0] = 1193ns;
slave_timing[0][192+20].t_rxd1[0][2] = 878ns;
slave_timing[0][192+20].t_rxd1[2][0] = 1479ns;
slave_timing[0][192+20].t_rxd2[0][2] = 1395ns;
slave_timing[0][192+20].t_rxd2[2][0] = 838ns;
slave_timing[0][192+20].t_rxd2[1][2] = 1087ns;
slave_timing[0][192+20].t_rxd2[2][1] = 1117ns;

slave_timing[0][192+21].info_corner          = 3;
slave_timing[0][192+21].info_temp__j__       = -40;
slave_timing[0][192+21].info_i__quite_rec__  = 0.000000000;
slave_timing[0][192+21].info_dtr__ib__       = -1;
slave_timing[0][192+21].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+21].info_i__max_slave__  = 0.025000000;
slave_timing[0][192+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][192+21].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+21].t_rxd1[0][1] = 1142ns;
slave_timing[0][192+21].t_rxd1[1][0] = 1230ns;
slave_timing[0][192+21].t_rxd1[0][2] = 854ns;
slave_timing[0][192+21].t_rxd1[2][0] = 1509ns;
slave_timing[0][192+21].t_rxd2[0][2] = 1296ns;
slave_timing[0][192+21].t_rxd2[2][0] = 892ns;
slave_timing[0][192+21].t_rxd2[1][2] = 964ns;
slave_timing[0][192+21].t_rxd2[2][1] = 1252ns;

slave_timing[0][192+22].info_corner          = 3;
slave_timing[0][192+22].info_temp__j__       = -40;
slave_timing[0][192+22].info_i__quite_rec__  = 0.000000000;
slave_timing[0][192+22].info_dtr__ib__       = 1;
slave_timing[0][192+22].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+22].info_i__max_slave__  = 0.023000000;
slave_timing[0][192+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][192+22].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+22].t_rxd1[0][1] = 1226ns;
slave_timing[0][192+22].t_rxd1[1][0] = 1155ns;
slave_timing[0][192+22].t_rxd1[0][2] = 891ns;
slave_timing[0][192+22].t_rxd1[2][0] = 1445ns;
slave_timing[0][192+22].t_rxd2[0][2] = 1488ns;
slave_timing[0][192+22].t_rxd2[2][0] = 786ns;
slave_timing[0][192+22].t_rxd2[1][2] = 1196ns;
slave_timing[0][192+22].t_rxd2[2][1] = 1021ns;

slave_timing[0][192+23].info_corner          = 3;
slave_timing[0][192+23].info_temp__j__       = -40;
slave_timing[0][192+23].info_i__quite_rec__  = 0.000000000;
slave_timing[0][192+23].info_dtr__ib__       = 1;
slave_timing[0][192+23].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+23].info_i__max_slave__  = 0.025000000;
slave_timing[0][192+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][192+23].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+23].t_rxd1[0][1] = 1169ns;
slave_timing[0][192+23].t_rxd1[1][0] = 1193ns;
slave_timing[0][192+23].t_rxd1[0][2] = 865ns;
slave_timing[0][192+23].t_rxd1[2][0] = 1477ns;
slave_timing[0][192+23].t_rxd2[0][2] = 1362ns;
slave_timing[0][192+23].t_rxd2[2][0] = 847ns;
slave_timing[0][192+23].t_rxd2[1][2] = 1051ns;
slave_timing[0][192+23].t_rxd2[2][1] = 1145ns;

slave_timing[0][192+24].info_corner          = 3;
slave_timing[0][192+24].info_temp__j__       = -40;
slave_timing[0][192+24].info_i__quite_rec__  = 0.040000000;
slave_timing[0][192+24].info_dtr__ib__       = -1;
slave_timing[0][192+24].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+24].info_i__max_slave__  = 0.023000000;
slave_timing[0][192+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][192+24].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+24].t_rxd1[0][1] = 1096ns;
slave_timing[0][192+24].t_rxd1[1][0] = 1098ns;
slave_timing[0][192+24].t_rxd1[0][2] = 805ns;
slave_timing[0][192+24].t_rxd1[2][0] = 1390ns;
slave_timing[0][192+24].t_rxd2[0][2] = 1364ns;
slave_timing[0][192+24].t_rxd2[2][0] = 815ns;
slave_timing[0][192+24].t_rxd2[1][2] = 1077ns;
slave_timing[0][192+24].t_rxd2[2][1] = 1102ns;

slave_timing[0][192+25].info_corner          = 3;
slave_timing[0][192+25].info_temp__j__       = -40;
slave_timing[0][192+25].info_i__quite_rec__  = 0.040000000;
slave_timing[0][192+25].info_dtr__ib__       = -1;
slave_timing[0][192+25].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+25].info_i__max_slave__  = 0.025000000;
slave_timing[0][192+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][192+25].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+25].t_rxd1[0][1] = 1048ns;
slave_timing[0][192+25].t_rxd1[1][0] = 1136ns;
slave_timing[0][192+25].t_rxd1[0][2] = 783ns;
slave_timing[0][192+25].t_rxd1[2][0] = 1422ns;
slave_timing[0][192+25].t_rxd2[0][2] = 1266ns;
slave_timing[0][192+25].t_rxd2[2][0] = 869ns;
slave_timing[0][192+25].t_rxd2[1][2] = 951ns;
slave_timing[0][192+25].t_rxd2[2][1] = 1235ns;

slave_timing[0][192+26].info_corner          = 3;
slave_timing[0][192+26].info_temp__j__       = -40;
slave_timing[0][192+26].info_i__quite_rec__  = 0.040000000;
slave_timing[0][192+26].info_dtr__ib__       = 1;
slave_timing[0][192+26].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+26].info_i__max_slave__  = 0.023000000;
slave_timing[0][192+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][192+26].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+26].t_rxd1[0][1] = 1130ns;
slave_timing[0][192+26].t_rxd1[1][0] = 1074ns;
slave_timing[0][192+26].t_rxd1[0][2] = 821ns;
slave_timing[0][192+26].t_rxd1[2][0] = 1370ns;
slave_timing[0][192+26].t_rxd2[0][2] = 1459ns;
slave_timing[0][192+26].t_rxd2[2][0] = 772ns;
slave_timing[0][192+26].t_rxd2[1][2] = 1183ns;
slave_timing[0][192+26].t_rxd2[2][1] = 1011ns;

slave_timing[0][192+27].info_corner          = 3;
slave_timing[0][192+27].info_temp__j__       = -40;
slave_timing[0][192+27].info_i__quite_rec__  = 0.040000000;
slave_timing[0][192+27].info_dtr__ib__       = 1;
slave_timing[0][192+27].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+27].info_i__max_slave__  = 0.025000000;
slave_timing[0][192+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[0][192+27].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+27].t_rxd1[0][1] = 1077ns;
slave_timing[0][192+27].t_rxd1[1][0] = 1109ns;
slave_timing[0][192+27].t_rxd1[0][2] = 798ns;
slave_timing[0][192+27].t_rxd1[2][0] = 1401ns;
slave_timing[0][192+27].t_rxd2[0][2] = 1334ns;
slave_timing[0][192+27].t_rxd2[2][0] = 831ns;
slave_timing[0][192+27].t_rxd2[1][2] = 1041ns;
slave_timing[0][192+27].t_rxd2[2][1] = 1139ns;

slave_timing[0][192+28].info_corner          = 3;
slave_timing[0][192+28].info_temp__j__       = -40;
slave_timing[0][192+28].info_i__quite_rec__  = 0.040000000;
slave_timing[0][192+28].info_dtr__ib__       = -1;
slave_timing[0][192+28].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+28].info_i__max_slave__  = 0.023000000;
slave_timing[0][192+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][192+28].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+28].t_rxd1[0][1] = 1140ns;
slave_timing[0][192+28].t_rxd1[1][0] = 1142ns;
slave_timing[0][192+28].t_rxd1[0][2] = 844ns;
slave_timing[0][192+28].t_rxd1[2][0] = 1429ns;
slave_timing[0][192+28].t_rxd2[0][2] = 1381ns;
slave_timing[0][192+28].t_rxd2[2][0] = 835ns;
slave_timing[0][192+28].t_rxd2[1][2] = 1091ns;
slave_timing[0][192+28].t_rxd2[2][1] = 1114ns;

slave_timing[0][192+29].info_corner          = 3;
slave_timing[0][192+29].info_temp__j__       = -40;
slave_timing[0][192+29].info_i__quite_rec__  = 0.040000000;
slave_timing[0][192+29].info_dtr__ib__       = -1;
slave_timing[0][192+29].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+29].info_i__max_slave__  = 0.025000000;
slave_timing[0][192+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][192+29].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+29].t_rxd1[0][1] = 1092ns;
slave_timing[0][192+29].t_rxd1[1][0] = 1178ns;
slave_timing[0][192+29].t_rxd1[0][2] = 809ns;
slave_timing[0][192+29].t_rxd1[2][0] = 1459ns;
slave_timing[0][192+29].t_rxd2[0][2] = 1269ns;
slave_timing[0][192+29].t_rxd2[2][0] = 888ns;
slave_timing[0][192+29].t_rxd2[1][2] = 973ns;
slave_timing[0][192+29].t_rxd2[2][1] = 1248ns;

slave_timing[0][192+30].info_corner          = 3;
slave_timing[0][192+30].info_temp__j__       = -40;
slave_timing[0][192+30].info_i__quite_rec__  = 0.040000000;
slave_timing[0][192+30].info_dtr__ib__       = 1;
slave_timing[0][192+30].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+30].info_i__max_slave__  = 0.023000000;
slave_timing[0][192+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][192+30].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+30].t_rxd1[0][1] = 1172ns;
slave_timing[0][192+30].t_rxd1[1][0] = 1115ns;
slave_timing[0][192+30].t_rxd1[0][2] = 857ns;
slave_timing[0][192+30].t_rxd1[2][0] = 1404ns;
slave_timing[0][192+30].t_rxd2[0][2] = 1474ns;
slave_timing[0][192+30].t_rxd2[2][0] = 788ns;
slave_timing[0][192+30].t_rxd2[1][2] = 1196ns;
slave_timing[0][192+30].t_rxd2[2][1] = 1020ns;

slave_timing[0][192+31].info_corner          = 3;
slave_timing[0][192+31].info_temp__j__       = -40;
slave_timing[0][192+31].info_i__quite_rec__  = 0.040000000;
slave_timing[0][192+31].info_dtr__ib__       = 1;
slave_timing[0][192+31].info_i__offset_rec__ = 0.000000000;
slave_timing[0][192+31].info_i__max_slave__  = 0.025000000;
slave_timing[0][192+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[0][192+31].info_r__dsi_bus__    = 5.000;

slave_timing[0][192+31].t_rxd1[0][1] = 1119ns;
slave_timing[0][192+31].t_rxd1[1][0] = 1152ns;
slave_timing[0][192+31].t_rxd1[0][2] = 832ns;
slave_timing[0][192+31].t_rxd1[2][0] = 1434ns;
slave_timing[0][192+31].t_rxd2[0][2] = 1349ns;
slave_timing[0][192+31].t_rxd2[2][0] = 848ns;
slave_timing[0][192+31].t_rxd2[1][2] = 1054ns;
slave_timing[0][192+31].t_rxd2[2][1] = 1147ns;


slave_timing[1][64+0].info_corner          = 3;
slave_timing[1][64+0].info_temp__j__       = 125;
slave_timing[1][64+0].info_i__quite_rec__  = 0.006000000;
slave_timing[1][64+0].info_dtr__ib__       = -1;
slave_timing[1][64+0].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+0].info_i__max_slave__  = 0.023000000;
slave_timing[1][64+0].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][64+0].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+0].t_rxd1[0][1] = 1653ns;
slave_timing[1][64+0].t_rxd1[1][0] = 1637ns;
slave_timing[1][64+0].t_rxd1[0][2] = 1236ns;
slave_timing[1][64+0].t_rxd1[2][0] = 1981ns;
slave_timing[1][64+0].t_rxd2[0][2] = 1965ns;
slave_timing[1][64+0].t_rxd2[2][0] = 1244ns;
slave_timing[1][64+0].t_rxd2[1][2] = 1652ns;
slave_timing[1][64+0].t_rxd2[2][1] = 1638ns;

slave_timing[1][64+1].info_corner          = 3;
slave_timing[1][64+1].info_temp__j__       = 125;
slave_timing[1][64+1].info_i__quite_rec__  = 0.006000000;
slave_timing[1][64+1].info_dtr__ib__       = -1;
slave_timing[1][64+1].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+1].info_i__max_slave__  = 0.025000000;
slave_timing[1][64+1].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][64+1].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+1].t_rxd1[0][1] = 1592ns;
slave_timing[1][64+1].t_rxd1[1][0] = 1685ns;
slave_timing[1][64+1].t_rxd1[0][2] = 1213ns;
slave_timing[1][64+1].t_rxd1[2][0] = 2014ns;
slave_timing[1][64+1].t_rxd2[0][2] = 1866ns;
slave_timing[1][64+1].t_rxd2[2][0] = 1326ns;
slave_timing[1][64+1].t_rxd2[1][2] = 1478ns;
slave_timing[1][64+1].t_rxd2[2][1] = 1805ns;

slave_timing[1][64+2].info_corner          = 3;
slave_timing[1][64+2].info_temp__j__       = 125;
slave_timing[1][64+2].info_i__quite_rec__  = 0.006000000;
slave_timing[1][64+2].info_dtr__ib__       = 1;
slave_timing[1][64+2].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+2].info_i__max_slave__  = 0.023000000;
slave_timing[1][64+2].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][64+2].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+2].t_rxd1[0][1] = 1679ns;
slave_timing[1][64+2].t_rxd1[1][0] = 1582ns;
slave_timing[1][64+2].t_rxd1[0][2] = 1255ns;
slave_timing[1][64+2].t_rxd1[2][0] = 1931ns;
slave_timing[1][64+2].t_rxd2[0][2] = 2071ns;
slave_timing[1][64+2].t_rxd2[2][0] = 1166ns;
slave_timing[1][64+2].t_rxd2[1][2] = 1789ns;
slave_timing[1][64+2].t_rxd2[2][1] = 1500ns;

slave_timing[1][64+3].info_corner          = 3;
slave_timing[1][64+3].info_temp__j__       = 125;
slave_timing[1][64+3].info_i__quite_rec__  = 0.006000000;
slave_timing[1][64+3].info_dtr__ib__       = 1;
slave_timing[1][64+3].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+3].info_i__max_slave__  = 0.025000000;
slave_timing[1][64+3].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][64+3].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+3].t_rxd1[0][1] = 1612ns;
slave_timing[1][64+3].t_rxd1[1][0] = 1631ns;
slave_timing[1][64+3].t_rxd1[0][2] = 1220ns;
slave_timing[1][64+3].t_rxd1[2][0] = 1963ns;
slave_timing[1][64+3].t_rxd2[0][2] = 1927ns;
slave_timing[1][64+3].t_rxd2[2][0] = 1256ns;
slave_timing[1][64+3].t_rxd2[1][2] = 1594ns;
slave_timing[1][64+3].t_rxd2[2][1] = 1663ns;

slave_timing[1][64+4].info_corner          = 3;
slave_timing[1][64+4].info_temp__j__       = 125;
slave_timing[1][64+4].info_i__quite_rec__  = 0.006000000;
slave_timing[1][64+4].info_dtr__ib__       = -1;
slave_timing[1][64+4].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+4].info_i__max_slave__  = 0.023000000;
slave_timing[1][64+4].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][64+4].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+4].t_rxd1[0][1] = 1858ns;
slave_timing[1][64+4].t_rxd1[1][0] = 1785ns;
slave_timing[1][64+4].t_rxd1[0][2] = 1408ns;
slave_timing[1][64+4].t_rxd1[2][0] = 2120ns;
slave_timing[1][64+4].t_rxd2[0][2] = 2033ns;
slave_timing[1][64+4].t_rxd2[2][0] = 1281ns;
slave_timing[1][64+4].t_rxd2[1][2] = 1681ns;
slave_timing[1][64+4].t_rxd2[2][1] = 1667ns;

slave_timing[1][64+5].info_corner          = 3;
slave_timing[1][64+5].info_temp__j__       = 125;
slave_timing[1][64+5].info_i__quite_rec__  = 0.006000000;
slave_timing[1][64+5].info_dtr__ib__       = -1;
slave_timing[1][64+5].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+5].info_i__max_slave__  = 0.025000000;
slave_timing[1][64+5].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][64+5].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+5].t_rxd1[0][1] = 1786ns;
slave_timing[1][64+5].t_rxd1[1][0] = 1829ns;
slave_timing[1][64+5].t_rxd1[0][2] = 1369ns;
slave_timing[1][64+5].t_rxd1[2][0] = 2151ns;
slave_timing[1][64+5].t_rxd2[0][2] = 1918ns;
slave_timing[1][64+5].t_rxd2[2][0] = 1359ns;
slave_timing[1][64+5].t_rxd2[1][2] = 1511ns;
slave_timing[1][64+5].t_rxd2[2][1] = 1831ns;

slave_timing[1][64+6].info_corner          = 3;
slave_timing[1][64+6].info_temp__j__       = 125;
slave_timing[1][64+6].info_i__quite_rec__  = 0.006000000;
slave_timing[1][64+6].info_dtr__ib__       = 1;
slave_timing[1][64+6].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+6].info_i__max_slave__  = 0.023000000;
slave_timing[1][64+6].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][64+6].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+6].t_rxd1[0][1] = 1874ns;
slave_timing[1][64+6].t_rxd1[1][0] = 1722ns;
slave_timing[1][64+6].t_rxd1[0][2] = 1407ns;
slave_timing[1][64+6].t_rxd1[2][0] = 2062ns;
slave_timing[1][64+6].t_rxd2[0][2] = 2113ns;
slave_timing[1][64+6].t_rxd2[2][0] = 1196ns;
slave_timing[1][64+6].t_rxd2[1][2] = 1811ns;
slave_timing[1][64+6].t_rxd2[2][1] = 1527ns;

slave_timing[1][64+7].info_corner          = 3;
slave_timing[1][64+7].info_temp__j__       = 125;
slave_timing[1][64+7].info_i__quite_rec__  = 0.006000000;
slave_timing[1][64+7].info_dtr__ib__       = 1;
slave_timing[1][64+7].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+7].info_i__max_slave__  = 0.025000000;
slave_timing[1][64+7].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][64+7].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+7].t_rxd1[0][1] = 1800ns;
slave_timing[1][64+7].t_rxd1[1][0] = 1769ns;
slave_timing[1][64+7].t_rxd1[0][2] = 1368ns;
slave_timing[1][64+7].t_rxd1[2][0] = 2093ns;
slave_timing[1][64+7].t_rxd2[0][2] = 1974ns;
slave_timing[1][64+7].t_rxd2[2][0] = 1289ns;
slave_timing[1][64+7].t_rxd2[1][2] = 1620ns;
slave_timing[1][64+7].t_rxd2[2][1] = 1690ns;

slave_timing[1][64+8].info_corner          = 3;
slave_timing[1][64+8].info_temp__j__       = 125;
slave_timing[1][64+8].info_i__quite_rec__  = 0.003000000;
slave_timing[1][64+8].info_dtr__ib__       = -1;
slave_timing[1][64+8].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+8].info_i__max_slave__  = 0.023000000;
slave_timing[1][64+8].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][64+8].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+8].t_rxd1[0][1] = 1606ns;
slave_timing[1][64+8].t_rxd1[1][0] = 1626ns;
slave_timing[1][64+8].t_rxd1[0][2] = 1215ns;
slave_timing[1][64+8].t_rxd1[2][0] = 1953ns;
slave_timing[1][64+8].t_rxd2[0][2] = 1940ns;
slave_timing[1][64+8].t_rxd2[2][0] = 1233ns;
slave_timing[1][64+8].t_rxd2[1][2] = 1619ns;
slave_timing[1][64+8].t_rxd2[2][1] = 1621ns;

slave_timing[1][64+9].info_corner          = 3;
slave_timing[1][64+9].info_temp__j__       = 125;
slave_timing[1][64+9].info_i__quite_rec__  = 0.003000000;
slave_timing[1][64+9].info_dtr__ib__       = -1;
slave_timing[1][64+9].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+9].info_i__max_slave__  = 0.025000000;
slave_timing[1][64+9].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][64+9].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+9].t_rxd1[0][1] = 1547ns;
slave_timing[1][64+9].t_rxd1[1][0] = 1670ns;
slave_timing[1][64+9].t_rxd1[0][2] = 1182ns;
slave_timing[1][64+9].t_rxd1[2][0] = 1983ns;
slave_timing[1][64+9].t_rxd2[0][2] = 1826ns;
slave_timing[1][64+9].t_rxd2[2][0] = 1311ns;
slave_timing[1][64+9].t_rxd2[1][2] = 1453ns;
slave_timing[1][64+9].t_rxd2[2][1] = 1783ns;

slave_timing[1][64+10].info_corner          = 3;
slave_timing[1][64+10].info_temp__j__       = 125;
slave_timing[1][64+10].info_i__quite_rec__  = 0.003000000;
slave_timing[1][64+10].info_dtr__ib__       = 1;
slave_timing[1][64+10].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+10].info_i__max_slave__  = 0.023000000;
slave_timing[1][64+10].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][64+10].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+10].t_rxd1[0][1] = 1653ns;
slave_timing[1][64+10].t_rxd1[1][0] = 1544ns;
slave_timing[1][64+10].t_rxd1[0][2] = 1234ns;
slave_timing[1][64+10].t_rxd1[2][0] = 1884ns;
slave_timing[1][64+10].t_rxd2[0][2] = 2042ns;
slave_timing[1][64+10].t_rxd2[2][0] = 1140ns;
slave_timing[1][64+10].t_rxd2[1][2] = 1776ns;
slave_timing[1][64+10].t_rxd2[2][1] = 1463ns;

slave_timing[1][64+11].info_corner          = 3;
slave_timing[1][64+11].info_temp__j__       = 125;
slave_timing[1][64+11].info_i__quite_rec__  = 0.003000000;
slave_timing[1][64+11].info_dtr__ib__       = 1;
slave_timing[1][64+11].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+11].info_i__max_slave__  = 0.025000000;
slave_timing[1][64+11].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][64+11].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+11].t_rxd1[0][1] = 1583ns;
slave_timing[1][64+11].t_rxd1[1][0] = 1590ns;
slave_timing[1][64+11].t_rxd1[0][2] = 1197ns;
slave_timing[1][64+11].t_rxd1[2][0] = 1916ns;
slave_timing[1][64+11].t_rxd2[0][2] = 1903ns;
slave_timing[1][64+11].t_rxd2[2][0] = 1231ns;
slave_timing[1][64+11].t_rxd2[1][2] = 1580ns;
slave_timing[1][64+11].t_rxd2[2][1] = 1625ns;

slave_timing[1][64+12].info_corner          = 3;
slave_timing[1][64+12].info_temp__j__       = 125;
slave_timing[1][64+12].info_i__quite_rec__  = 0.003000000;
slave_timing[1][64+12].info_dtr__ib__       = -1;
slave_timing[1][64+12].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+12].info_i__max_slave__  = 0.023000000;
slave_timing[1][64+12].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][64+12].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+12].t_rxd1[0][1] = 1822ns;
slave_timing[1][64+12].t_rxd1[1][0] = 1774ns;
slave_timing[1][64+12].t_rxd1[0][2] = 1387ns;
slave_timing[1][64+12].t_rxd1[2][0] = 2092ns;
slave_timing[1][64+12].t_rxd2[0][2] = 1985ns;
slave_timing[1][64+12].t_rxd2[2][0] = 1265ns;
slave_timing[1][64+12].t_rxd2[1][2] = 1669ns;
slave_timing[1][64+12].t_rxd2[2][1] = 1626ns;

slave_timing[1][64+13].info_corner          = 3;
slave_timing[1][64+13].info_temp__j__       = 125;
slave_timing[1][64+13].info_i__quite_rec__  = 0.003000000;
slave_timing[1][64+13].info_dtr__ib__       = -1;
slave_timing[1][64+13].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+13].info_i__max_slave__  = 0.025000000;
slave_timing[1][64+13].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][64+13].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+13].t_rxd1[0][1] = 1752ns;
slave_timing[1][64+13].t_rxd1[1][0] = 1817ns;
slave_timing[1][64+13].t_rxd1[0][2] = 1349ns;
slave_timing[1][64+13].t_rxd1[2][0] = 2121ns;
slave_timing[1][64+13].t_rxd2[0][2] = 1875ns;
slave_timing[1][64+13].t_rxd2[2][0] = 1344ns;
slave_timing[1][64+13].t_rxd2[1][2] = 1502ns;
slave_timing[1][64+13].t_rxd2[2][1] = 1788ns;

slave_timing[1][64+14].info_corner          = 3;
slave_timing[1][64+14].info_temp__j__       = 125;
slave_timing[1][64+14].info_i__quite_rec__  = 0.003000000;
slave_timing[1][64+14].info_dtr__ib__       = 1;
slave_timing[1][64+14].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+14].info_i__max_slave__  = 0.023000000;
slave_timing[1][64+14].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][64+14].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+14].t_rxd1[0][1] = 1861ns;
slave_timing[1][64+14].t_rxd1[1][0] = 1681ns;
slave_timing[1][64+14].t_rxd1[0][2] = 1400ns;
slave_timing[1][64+14].t_rxd1[2][0] = 2013ns;
slave_timing[1][64+14].t_rxd2[0][2] = 2080ns;
slave_timing[1][64+14].t_rxd2[2][0] = 1172ns;
slave_timing[1][64+14].t_rxd2[1][2] = 1796ns;
slave_timing[1][64+14].t_rxd2[2][1] = 1490ns;

slave_timing[1][64+15].info_corner          = 3;
slave_timing[1][64+15].info_temp__j__       = 125;
slave_timing[1][64+15].info_i__quite_rec__  = 0.003000000;
slave_timing[1][64+15].info_dtr__ib__       = 1;
slave_timing[1][64+15].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+15].info_i__max_slave__  = 0.025000000;
slave_timing[1][64+15].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][64+15].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+15].t_rxd1[0][1] = 1790ns;
slave_timing[1][64+15].t_rxd1[1][0] = 1729ns;
slave_timing[1][64+15].t_rxd1[0][2] = 1361ns;
slave_timing[1][64+15].t_rxd1[2][0] = 2045ns;
slave_timing[1][64+15].t_rxd2[0][2] = 1944ns;
slave_timing[1][64+15].t_rxd2[2][0] = 1260ns;
slave_timing[1][64+15].t_rxd2[1][2] = 1607ns;
slave_timing[1][64+15].t_rxd2[2][1] = 1644ns;

slave_timing[1][64+16].info_corner          = 3;
slave_timing[1][64+16].info_temp__j__       = 125;
slave_timing[1][64+16].info_i__quite_rec__  = 0.000000000;
slave_timing[1][64+16].info_dtr__ib__       = -1;
slave_timing[1][64+16].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+16].info_i__max_slave__  = 0.023000000;
slave_timing[1][64+16].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][64+16].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+16].t_rxd1[0][1] = 1588ns;
slave_timing[1][64+16].t_rxd1[1][0] = 1585ns;
slave_timing[1][64+16].t_rxd1[0][2] = 1199ns;
slave_timing[1][64+16].t_rxd1[2][0] = 1897ns;
slave_timing[1][64+16].t_rxd2[0][2] = 1903ns;
slave_timing[1][64+16].t_rxd2[2][0] = 1207ns;
slave_timing[1][64+16].t_rxd2[1][2] = 1599ns;
slave_timing[1][64+16].t_rxd2[2][1] = 1585ns;

slave_timing[1][64+17].info_corner          = 3;
slave_timing[1][64+17].info_temp__j__       = 125;
slave_timing[1][64+17].info_i__quite_rec__  = 0.000000000;
slave_timing[1][64+17].info_dtr__ib__       = -1;
slave_timing[1][64+17].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+17].info_i__max_slave__  = 0.025000000;
slave_timing[1][64+17].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][64+17].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+17].t_rxd1[0][1] = 1528ns;
slave_timing[1][64+17].t_rxd1[1][0] = 1626ns;
slave_timing[1][64+17].t_rxd1[0][2] = 1166ns;
slave_timing[1][64+17].t_rxd1[2][0] = 1929ns;
slave_timing[1][64+17].t_rxd2[0][2] = 1793ns;
slave_timing[1][64+17].t_rxd2[2][0] = 1286ns;
slave_timing[1][64+17].t_rxd2[1][2] = 1434ns;
slave_timing[1][64+17].t_rxd2[2][1] = 1745ns;

slave_timing[1][64+18].info_corner          = 3;
slave_timing[1][64+18].info_temp__j__       = 125;
slave_timing[1][64+18].info_i__quite_rec__  = 0.000000000;
slave_timing[1][64+18].info_dtr__ib__       = 1;
slave_timing[1][64+18].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+18].info_i__max_slave__  = 0.023000000;
slave_timing[1][64+18].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][64+18].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+18].t_rxd1[0][1] = 1637ns;
slave_timing[1][64+18].t_rxd1[1][0] = 1510ns;
slave_timing[1][64+18].t_rxd1[0][2] = 1219ns;
slave_timing[1][64+18].t_rxd1[2][0] = 1837ns;
slave_timing[1][64+18].t_rxd2[0][2] = 2005ns;
slave_timing[1][64+18].t_rxd2[2][0] = 1112ns;
slave_timing[1][64+18].t_rxd2[1][2] = 1747ns;
slave_timing[1][64+18].t_rxd2[2][1] = 1427ns;

slave_timing[1][64+19].info_corner          = 3;
slave_timing[1][64+19].info_temp__j__       = 125;
slave_timing[1][64+19].info_i__quite_rec__  = 0.000000000;
slave_timing[1][64+19].info_dtr__ib__       = 1;
slave_timing[1][64+19].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+19].info_i__max_slave__  = 0.025000000;
slave_timing[1][64+19].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][64+19].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+19].t_rxd1[0][1] = 1569ns;
slave_timing[1][64+19].t_rxd1[1][0] = 1553ns;
slave_timing[1][64+19].t_rxd1[0][2] = 1182ns;
slave_timing[1][64+19].t_rxd1[2][0] = 1868ns;
slave_timing[1][64+19].t_rxd2[0][2] = 1865ns;
slave_timing[1][64+19].t_rxd2[2][0] = 1204ns;
slave_timing[1][64+19].t_rxd2[1][2] = 1556ns;
slave_timing[1][64+19].t_rxd2[2][1] = 1585ns;

slave_timing[1][64+20].info_corner          = 3;
slave_timing[1][64+20].info_temp__j__       = 125;
slave_timing[1][64+20].info_i__quite_rec__  = 0.000000000;
slave_timing[1][64+20].info_dtr__ib__       = -1;
slave_timing[1][64+20].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+20].info_i__max_slave__  = 0.023000000;
slave_timing[1][64+20].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][64+20].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+20].t_rxd1[0][1] = 1827ns;
slave_timing[1][64+20].t_rxd1[1][0] = 1727ns;
slave_timing[1][64+20].t_rxd1[0][2] = 1386ns;
slave_timing[1][64+20].t_rxd1[2][0] = 2029ns;
slave_timing[1][64+20].t_rxd2[0][2] = 1945ns;
slave_timing[1][64+20].t_rxd2[2][0] = 1238ns;
slave_timing[1][64+20].t_rxd2[1][2] = 1622ns;
slave_timing[1][64+20].t_rxd2[2][1] = 1609ns;

slave_timing[1][64+21].info_corner          = 3;
slave_timing[1][64+21].info_temp__j__       = 125;
slave_timing[1][64+21].info_i__quite_rec__  = 0.000000000;
slave_timing[1][64+21].info_dtr__ib__       = -1;
slave_timing[1][64+21].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+21].info_i__max_slave__  = 0.025000000;
slave_timing[1][64+21].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][64+21].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+21].t_rxd1[0][1] = 1758ns;
slave_timing[1][64+21].t_rxd1[1][0] = 1769ns;
slave_timing[1][64+21].t_rxd1[0][2] = 1348ns;
slave_timing[1][64+21].t_rxd1[2][0] = 2058ns;
slave_timing[1][64+21].t_rxd2[0][2] = 1837ns;
slave_timing[1][64+21].t_rxd2[2][0] = 1315ns;
slave_timing[1][64+21].t_rxd2[1][2] = 1460ns;
slave_timing[1][64+21].t_rxd2[2][1] = 1764ns;

slave_timing[1][64+22].info_corner          = 3;
slave_timing[1][64+22].info_temp__j__       = 125;
slave_timing[1][64+22].info_i__quite_rec__  = 0.000000000;
slave_timing[1][64+22].info_dtr__ib__       = 1;
slave_timing[1][64+22].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+22].info_i__max_slave__  = 0.023000000;
slave_timing[1][64+22].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][64+22].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+22].t_rxd1[0][1] = 1869ns;
slave_timing[1][64+22].t_rxd1[1][0] = 1647ns;
slave_timing[1][64+22].t_rxd1[0][2] = 1403ns;
slave_timing[1][64+22].t_rxd1[2][0] = 1963ns;
slave_timing[1][64+22].t_rxd2[0][2] = 2034ns;
slave_timing[1][64+22].t_rxd2[2][0] = 1142ns;
slave_timing[1][64+22].t_rxd2[1][2] = 1766ns;
slave_timing[1][64+22].t_rxd2[2][1] = 1453ns;

slave_timing[1][64+23].info_corner          = 3;
slave_timing[1][64+23].info_temp__j__       = 125;
slave_timing[1][64+23].info_i__quite_rec__  = 0.000000000;
slave_timing[1][64+23].info_dtr__ib__       = 1;
slave_timing[1][64+23].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+23].info_i__max_slave__  = 0.025000000;
slave_timing[1][64+23].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][64+23].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+23].t_rxd1[0][1] = 1795ns;
slave_timing[1][64+23].t_rxd1[1][0] = 1692ns;
slave_timing[1][64+23].t_rxd1[0][2] = 1364ns;
slave_timing[1][64+23].t_rxd1[2][0] = 1992ns;
slave_timing[1][64+23].t_rxd2[0][2] = 1902ns;
slave_timing[1][64+23].t_rxd2[2][0] = 1233ns;
slave_timing[1][64+23].t_rxd2[1][2] = 1581ns;
slave_timing[1][64+23].t_rxd2[2][1] = 1608ns;

slave_timing[1][64+24].info_corner          = 3;
slave_timing[1][64+24].info_temp__j__       = 125;
slave_timing[1][64+24].info_i__quite_rec__  = 0.040000000;
slave_timing[1][64+24].info_dtr__ib__       = -1;
slave_timing[1][64+24].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+24].info_i__max_slave__  = 0.023000000;
slave_timing[1][64+24].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][64+24].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+24].t_rxd1[0][1] = 1676ns;
slave_timing[1][64+24].t_rxd1[1][0] = 1680ns;
slave_timing[1][64+24].t_rxd1[0][2] = 1265ns;
slave_timing[1][64+24].t_rxd1[2][0] = 2019ns;
slave_timing[1][64+24].t_rxd2[0][2] = 2029ns;
slave_timing[1][64+24].t_rxd2[2][0] = 1277ns;
slave_timing[1][64+24].t_rxd2[1][2] = 1667ns;
slave_timing[1][64+24].t_rxd2[2][1] = 1654ns;

slave_timing[1][64+25].info_corner          = 3;
slave_timing[1][64+25].info_temp__j__       = 125;
slave_timing[1][64+25].info_i__quite_rec__  = 0.040000000;
slave_timing[1][64+25].info_dtr__ib__       = -1;
slave_timing[1][64+25].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+25].info_i__max_slave__  = 0.025000000;
slave_timing[1][64+25].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][64+25].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+25].t_rxd1[0][1] = 1611ns;
slave_timing[1][64+25].t_rxd1[1][0] = 1726ns;
slave_timing[1][64+25].t_rxd1[0][2] = 1231ns;
slave_timing[1][64+25].t_rxd1[2][0] = 2051ns;
slave_timing[1][64+25].t_rxd2[0][2] = 1922ns;
slave_timing[1][64+25].t_rxd2[2][0] = 1365ns;
slave_timing[1][64+25].t_rxd2[1][2] = 1500ns;
slave_timing[1][64+25].t_rxd2[2][1] = 1826ns;

slave_timing[1][64+26].info_corner          = 3;
slave_timing[1][64+26].info_temp__j__       = 125;
slave_timing[1][64+26].info_i__quite_rec__  = 0.040000000;
slave_timing[1][64+26].info_dtr__ib__       = 1;
slave_timing[1][64+26].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+26].info_i__max_slave__  = 0.023000000;
slave_timing[1][64+26].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][64+26].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+26].t_rxd1[0][1] = 1721ns;
slave_timing[1][64+26].t_rxd1[1][0] = 1642ns;
slave_timing[1][64+26].t_rxd1[0][2] = 1289ns;
slave_timing[1][64+26].t_rxd1[2][0] = 1991ns;
slave_timing[1][64+26].t_rxd2[0][2] = 2139ns;
slave_timing[1][64+26].t_rxd2[2][0] = 1211ns;
slave_timing[1][64+26].t_rxd2[1][2] = 1816ns;
slave_timing[1][64+26].t_rxd2[2][1] = 1538ns;

slave_timing[1][64+27].info_corner          = 3;
slave_timing[1][64+27].info_temp__j__       = 125;
slave_timing[1][64+27].info_i__quite_rec__  = 0.040000000;
slave_timing[1][64+27].info_dtr__ib__       = 1;
slave_timing[1][64+27].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+27].info_i__max_slave__  = 0.025000000;
slave_timing[1][64+27].info_c__dsi_bus__    = 0.000000010000;
slave_timing[1][64+27].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+27].t_rxd1[0][1] = 1652ns;
slave_timing[1][64+27].t_rxd1[1][0] = 1690ns;
slave_timing[1][64+27].t_rxd1[0][2] = 1253ns;
slave_timing[1][64+27].t_rxd1[2][0] = 2024ns;
slave_timing[1][64+27].t_rxd2[0][2] = 2007ns;
slave_timing[1][64+27].t_rxd2[2][0] = 1308ns;
slave_timing[1][64+27].t_rxd2[1][2] = 1629ns;
slave_timing[1][64+27].t_rxd2[2][1] = 1712ns;

slave_timing[1][64+28].info_corner          = 3;
slave_timing[1][64+28].info_temp__j__       = 125;
slave_timing[1][64+28].info_i__quite_rec__  = 0.040000000;
slave_timing[1][64+28].info_dtr__ib__       = -1;
slave_timing[1][64+28].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+28].info_i__max_slave__  = 0.023000000;
slave_timing[1][64+28].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][64+28].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+28].t_rxd1[0][1] = 1774ns;
slave_timing[1][64+28].t_rxd1[1][0] = 1761ns;
slave_timing[1][64+28].t_rxd1[0][2] = 1358ns;
slave_timing[1][64+28].t_rxd1[2][0] = 1984ns;
slave_timing[1][64+28].t_rxd2[0][2] = 2112ns;
slave_timing[1][64+28].t_rxd2[2][0] = 1577ns;
slave_timing[1][64+28].t_rxd2[1][2] = 1744ns;
slave_timing[1][64+28].t_rxd2[2][1] = 2002ns;

slave_timing[1][64+29].info_corner          = 3;
slave_timing[1][64+29].info_temp__j__       = 125;
slave_timing[1][64+29].info_i__quite_rec__  = 0.040000000;
slave_timing[1][64+29].info_dtr__ib__       = -1;
slave_timing[1][64+29].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+29].info_i__max_slave__  = 0.025000000;
slave_timing[1][64+29].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][64+29].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+29].t_rxd1[0][1] = 1709ns;
slave_timing[1][64+29].t_rxd1[1][0] = 1808ns;
slave_timing[1][64+29].t_rxd1[0][2] = 1322ns;
slave_timing[1][64+29].t_rxd1[2][0] = 2064ns;
slave_timing[1][64+29].t_rxd2[0][2] = 2018ns;
slave_timing[1][64+29].t_rxd2[2][0] = 1710ns;
slave_timing[1][64+29].t_rxd2[1][2] = 1582ns;
slave_timing[1][64+29].t_rxd2[2][1] = 2259ns;

slave_timing[1][64+30].info_corner          = 3;
slave_timing[1][64+30].info_temp__j__       = 125;
slave_timing[1][64+30].info_i__quite_rec__  = 0.040000000;
slave_timing[1][64+30].info_dtr__ib__       = 1;
slave_timing[1][64+30].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+30].info_i__max_slave__  = 0.023000000;
slave_timing[1][64+30].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][64+30].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+30].t_rxd1[0][1] = 1814ns;
slave_timing[1][64+30].t_rxd1[1][0] = 1719ns;
slave_timing[1][64+30].t_rxd1[0][2] = 1378ns;
slave_timing[1][64+30].t_rxd1[2][0] = 1956ns;
slave_timing[1][64+30].t_rxd2[0][2] = 2222ns;
slave_timing[1][64+30].t_rxd2[2][0] = 1488ns;
slave_timing[1][64+30].t_rxd2[1][2] = 1893ns;
slave_timing[1][64+30].t_rxd2[2][1] = 1860ns;

slave_timing[1][64+31].info_corner          = 3;
slave_timing[1][64+31].info_temp__j__       = 125;
slave_timing[1][64+31].info_i__quite_rec__  = 0.040000000;
slave_timing[1][64+31].info_dtr__ib__       = 1;
slave_timing[1][64+31].info_i__offset_rec__ = 0.000000000;
slave_timing[1][64+31].info_i__max_slave__  = 0.025000000;
slave_timing[1][64+31].info_c__dsi_bus__    = 0.000000050000;
slave_timing[1][64+31].info_r__dsi_bus__    = 5.000;

slave_timing[1][64+31].t_rxd1[0][1] = 1745ns;
slave_timing[1][64+31].t_rxd1[1][0] = 1767ns;
slave_timing[1][64+31].t_rxd1[0][2] = 1340ns;
slave_timing[1][64+31].t_rxd1[2][0] = 2024ns;
slave_timing[1][64+31].t_rxd2[0][2] = 2108ns;
slave_timing[1][64+31].t_rxd2[2][0] = 1629ns;
slave_timing[1][64+31].t_rxd2[1][2] = 1715ns;
slave_timing[1][64+31].t_rxd2[2][1] = 2111ns;
